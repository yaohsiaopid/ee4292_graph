module top
#(
    parameter K = 16,
    parameter D = 256,
    parameter DIST_BW = 1,
    parameter DIST_ADDR_SPACE = 16,
    parameter LOC_BW = 5,
    parameter LOC_ADDR_SPACE = 4,
    parameter NEXT_BW = 4,
    parameter NEXT_ADDR_SPACE = 4,
    parameter PRO_BW = 8,
    parameter PRO_ADDR_SPACE = 4,
    parameter VID_BW = 16,  
    parameter VID_ADDR_SPACE = 5,
    parameter Q = 16
)
(
    input clk, 
	input en,
    input rst_n,
	
	// K * vid_sram
	input [Q*VID_BW-1:0] vid_sram_rdata0, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr0,
	input [Q*VID_BW-1:0] vid_sram_rdata1, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr1,
	input [Q*VID_BW-1:0] vid_sram_rdata2, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr2,
	input [Q*VID_BW-1:0] vid_sram_rdata3, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr3,
	input [Q*VID_BW-1:0] vid_sram_rdata4, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr4,
	input [Q*VID_BW-1:0] vid_sram_rdata5, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr5,
	input [Q*VID_BW-1:0] vid_sram_rdata6, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr6,
	input [Q*VID_BW-1:0] vid_sram_rdata7, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr7,
	input [Q*VID_BW-1:0] vid_sram_rdata8, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr8,
	input [Q*VID_BW-1:0] vid_sram_rdata9, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr9,
	input [Q*VID_BW-1:0] vid_sram_rdata10, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr10,
	input [Q*VID_BW-1:0] vid_sram_rdata11, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr11,
	input [Q*VID_BW-1:0] vid_sram_rdata12, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr12,
	input [Q*VID_BW-1:0] vid_sram_rdata13, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr13,
	input [Q*VID_BW-1:0] vid_sram_rdata14, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr14,
	input [Q*VID_BW-1:0] vid_sram_rdata15, output reg [VID_ADDR_SPACE-1:0] vid_sram_raddr15,
	
	output [K-1:0] vidsram_wen,
	output [Q*VID_BW-1:0] vid_sram_wdata0, 	output [VID_ADDR_SPACE-1:0] vid_sram_waddr0,
	output [Q*VID_BW-1:0] vid_sram_wdata1, 	output [VID_ADDR_SPACE-1:0] vid_sram_waddr1,
	output [Q*VID_BW-1:0] vid_sram_wdata2, 	output [VID_ADDR_SPACE-1:0] vid_sram_waddr2,
	output [Q*VID_BW-1:0] vid_sram_wdata3, 	output [VID_ADDR_SPACE-1:0] vid_sram_waddr3,
	output [Q*VID_BW-1:0] vid_sram_wdata4, 	output [VID_ADDR_SPACE-1:0] vid_sram_waddr4,
	output [Q*VID_BW-1:0] vid_sram_wdata5, 	output [VID_ADDR_SPACE-1:0] vid_sram_waddr5,
	output [Q*VID_BW-1:0] vid_sram_wdata6, 	output [VID_ADDR_SPACE-1:0] vid_sram_waddr6,
	output [Q*VID_BW-1:0] vid_sram_wdata7, 	output [VID_ADDR_SPACE-1:0] vid_sram_waddr7,
	output [Q*VID_BW-1:0] vid_sram_wdata8, 	output [VID_ADDR_SPACE-1:0] vid_sram_waddr8,
	output [Q*VID_BW-1:0] vid_sram_wdata9, 	output [VID_ADDR_SPACE-1:0] vid_sram_waddr9,
	output [Q*VID_BW-1:0] vid_sram_wdata10, output [VID_ADDR_SPACE-1:0] vid_sram_waddr10,
	output [Q*VID_BW-1:0] vid_sram_wdata11, output [VID_ADDR_SPACE-1:0] vid_sram_waddr11,
	output [Q*VID_BW-1:0] vid_sram_wdata12, output [VID_ADDR_SPACE-1:0] vid_sram_waddr12,
	output [Q*VID_BW-1:0] vid_sram_wdata13, output [VID_ADDR_SPACE-1:0] vid_sram_waddr13,
	output [Q*VID_BW-1:0] vid_sram_wdata14, output [VID_ADDR_SPACE-1:0] vid_sram_waddr14,
	output [Q*VID_BW-1:0] vid_sram_wdata15, output [VID_ADDR_SPACE-1:0] vid_sram_waddr15,

	// K * loc_sram
	output reg loc_sram_wen,
	input [D*LOC_BW-1:0] loc_sram_rdata0, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr0,
	input [D*LOC_BW-1:0] loc_sram_rdata1, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr1,
	input [D*LOC_BW-1:0] loc_sram_rdata2, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr2,
	input [D*LOC_BW-1:0] loc_sram_rdata3, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr3,
	input [D*LOC_BW-1:0] loc_sram_rdata4, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr4,
	input [D*LOC_BW-1:0] loc_sram_rdata5, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr5,
	input [D*LOC_BW-1:0] loc_sram_rdata6, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr6,
	input [D*LOC_BW-1:0] loc_sram_rdata7, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr7,
	input [D*LOC_BW-1:0] loc_sram_rdata8, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr8,
	input [D*LOC_BW-1:0] loc_sram_rdata9, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr9,
	input [D*LOC_BW-1:0] loc_sram_rdata10, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr10,
	input [D*LOC_BW-1:0] loc_sram_rdata11, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr11,
	input [D*LOC_BW-1:0] loc_sram_rdata12, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr12,
	input [D*LOC_BW-1:0] loc_sram_rdata13, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr13,
	input [D*LOC_BW-1:0] loc_sram_rdata14, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr14,
	input [D*LOC_BW-1:0] loc_sram_rdata15, output [LOC_ADDR_SPACE-1:0] loc_sram_raddr15,

	
	output reg [D*LOC_BW-1:0] loc_sram_wdata0, 	output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr0, output reg [D-1:0] loc_wbytemask0,
	output reg [D*LOC_BW-1:0] loc_sram_wdata1, 	output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr1, output reg [D-1:0] loc_wbytemask1,
	output reg [D*LOC_BW-1:0] loc_sram_wdata2, 	output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr2, output reg [D-1:0] loc_wbytemask2,
	output reg [D*LOC_BW-1:0] loc_sram_wdata3, 	output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr3, output reg [D-1:0] loc_wbytemask3,
	output reg [D*LOC_BW-1:0] loc_sram_wdata4, 	output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr4, output reg [D-1:0] loc_wbytemask4,
	output reg [D*LOC_BW-1:0] loc_sram_wdata5, 	output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr5, output reg [D-1:0] loc_wbytemask5,
	output reg [D*LOC_BW-1:0] loc_sram_wdata6, 	output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr6, output reg [D-1:0] loc_wbytemask6,
	output reg [D*LOC_BW-1:0] loc_sram_wdata7, 	output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr7, output reg [D-1:0] loc_wbytemask7,
	output reg [D*LOC_BW-1:0] loc_sram_wdata8, 	output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr8, output reg [D-1:0] loc_wbytemask8,
	output reg [D*LOC_BW-1:0] loc_sram_wdata9, 	output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr9, output reg [D-1:0] loc_wbytemask9,
	output reg [D*LOC_BW-1:0] loc_sram_wdata10, output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr10, output reg [D-1:0] loc_wbytemask10,
	output reg [D*LOC_BW-1:0] loc_sram_wdata11, output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr11, output reg [D-1:0] loc_wbytemask11,
	output reg [D*LOC_BW-1:0] loc_sram_wdata12, output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr12, output reg [D-1:0] loc_wbytemask12,
	output reg [D*LOC_BW-1:0] loc_sram_wdata13, output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr13, output reg [D-1:0] loc_wbytemask13,
	output reg [D*LOC_BW-1:0] loc_sram_wdata14, output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr14, output reg [D-1:0] loc_wbytemask14,
	output reg [D*LOC_BW-1:0] loc_sram_wdata15, output reg [LOC_ADDR_SPACE-1:0] loc_sram_waddr15, output reg [D-1:0] loc_wbytemask15,

	// K * dist_sram
	input [D*DIST_BW-1:0] dist_sram_rdata0, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr0,
	input [D*DIST_BW-1:0] dist_sram_rdata1, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr1,
	input [D*DIST_BW-1:0] dist_sram_rdata2, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr2,
	input [D*DIST_BW-1:0] dist_sram_rdata3, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr3,
	input [D*DIST_BW-1:0] dist_sram_rdata4, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr4,
	input [D*DIST_BW-1:0] dist_sram_rdata5, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr5,
	input [D*DIST_BW-1:0] dist_sram_rdata6, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr6,
	input [D*DIST_BW-1:0] dist_sram_rdata7, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr7,
	input [D*DIST_BW-1:0] dist_sram_rdata8, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr8,
	input [D*DIST_BW-1:0] dist_sram_rdata9, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr9,
	input [D*DIST_BW-1:0] dist_sram_rdata10, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr10,
	input [D*DIST_BW-1:0] dist_sram_rdata11, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr11,
	input [D*DIST_BW-1:0] dist_sram_rdata12, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr12,
	input [D*DIST_BW-1:0] dist_sram_rdata13, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr13,
	input [D*DIST_BW-1:0] dist_sram_rdata14, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr14,
	input [D*DIST_BW-1:0] dist_sram_rdata15, output [DIST_ADDR_SPACE-1:0] dist_sram_raddr15,

	// K * next_sram
	output worker_wen,
	input [Q*NEXT_BW-1:0] next_sram_rdata0, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr0,
	input [Q*NEXT_BW-1:0] next_sram_rdata1, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr1,
	input [Q*NEXT_BW-1:0] next_sram_rdata2, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr2,
	input [Q*NEXT_BW-1:0] next_sram_rdata3, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr3,
	input [Q*NEXT_BW-1:0] next_sram_rdata4, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr4,
	input [Q*NEXT_BW-1:0] next_sram_rdata5, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr5,
	input [Q*NEXT_BW-1:0] next_sram_rdata6, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr6,
	input [Q*NEXT_BW-1:0] next_sram_rdata7, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr7,
	input [Q*NEXT_BW-1:0] next_sram_rdata8, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr8,
	input [Q*NEXT_BW-1:0] next_sram_rdata9, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr9,
	input [Q*NEXT_BW-1:0] next_sram_rdata10, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr10,
	input [Q*NEXT_BW-1:0] next_sram_rdata11, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr11,
	input [Q*NEXT_BW-1:0] next_sram_rdata12, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr12,
	input [Q*NEXT_BW-1:0] next_sram_rdata13, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr13,
	input [Q*NEXT_BW-1:0] next_sram_rdata14, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr14,
	input [Q*NEXT_BW-1:0] next_sram_rdata15, output [NEXT_ADDR_SPACE-1:0] next_sram_raddr15,

	output [Q*NEXT_BW-1:0] next_sram_wdata0, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr0, output [Q-1:0] next_wbytemask0,
	output [Q*NEXT_BW-1:0] next_sram_wdata1, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr1, output [Q-1:0] next_wbytemask1,
	output [Q*NEXT_BW-1:0] next_sram_wdata2, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr2, output [Q-1:0] next_wbytemask2,
	output [Q*NEXT_BW-1:0] next_sram_wdata3, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr3, output [Q-1:0] next_wbytemask3,
	output [Q*NEXT_BW-1:0] next_sram_wdata4, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr4, output [Q-1:0] next_wbytemask4,
	output [Q*NEXT_BW-1:0] next_sram_wdata5, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr5, output [Q-1:0] next_wbytemask5,
	output [Q*NEXT_BW-1:0] next_sram_wdata6, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr6, output [Q-1:0] next_wbytemask6,
	output [Q*NEXT_BW-1:0] next_sram_wdata7, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr7, output [Q-1:0] next_wbytemask7,
	output [Q*NEXT_BW-1:0] next_sram_wdata8, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr8, output [Q-1:0] next_wbytemask8,
	output [Q*NEXT_BW-1:0] next_sram_wdata9, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr9, output [Q-1:0] next_wbytemask9,
	output [Q*NEXT_BW-1:0] next_sram_wdata10, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr10, output [Q-1:0] next_wbytemask10,
	output [Q*NEXT_BW-1:0] next_sram_wdata11, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr11, output [Q-1:0] next_wbytemask11,
	output [Q*NEXT_BW-1:0] next_sram_wdata12, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr12, output [Q-1:0] next_wbytemask12,
	output [Q*NEXT_BW-1:0] next_sram_wdata13, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr13, output [Q-1:0] next_wbytemask13,
	output [Q*NEXT_BW-1:0] next_sram_wdata14, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr14, output [Q-1:0] next_wbytemask14,
	output [Q*NEXT_BW-1:0] next_sram_wdata15, output [NEXT_ADDR_SPACE-1:0] next_sram_waddr15, output [Q-1:0] next_wbytemask15,

	// K * pro_sram
	input [Q*PRO_BW-1:0] pro_sram_rdata0, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr0,
	input [Q*PRO_BW-1:0] pro_sram_rdata1, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr1,
	input [Q*PRO_BW-1:0] pro_sram_rdata2, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr2,
	input [Q*PRO_BW-1:0] pro_sram_rdata3, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr3,
	input [Q*PRO_BW-1:0] pro_sram_rdata4, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr4,
	input [Q*PRO_BW-1:0] pro_sram_rdata5, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr5,
	input [Q*PRO_BW-1:0] pro_sram_rdata6, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr6,
	input [Q*PRO_BW-1:0] pro_sram_rdata7, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr7,
	input [Q*PRO_BW-1:0] pro_sram_rdata8, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr8,
	input [Q*PRO_BW-1:0] pro_sram_rdata9, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr9,
	input [Q*PRO_BW-1:0] pro_sram_rdata10, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr10,
	input [Q*PRO_BW-1:0] pro_sram_rdata11, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr11,
	input [Q*PRO_BW-1:0] pro_sram_rdata12, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr12,
	input [Q*PRO_BW-1:0] pro_sram_rdata13, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr13,
	input [Q*PRO_BW-1:0] pro_sram_rdata14, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr14,
	input [Q*PRO_BW-1:0] pro_sram_rdata15, output [PRO_ADDR_SPACE-1:0] pro_sram_raddr15,

	output [Q*PRO_BW-1:0] pro_sram_wdata0, 	output [PRO_ADDR_SPACE-1:0] pro_sram_waddr0, output [Q-1:0] pro_wbytemask0,
	output [Q*PRO_BW-1:0] pro_sram_wdata1, 	output [PRO_ADDR_SPACE-1:0] pro_sram_waddr1, output [Q-1:0] pro_wbytemask1,
	output [Q*PRO_BW-1:0] pro_sram_wdata2, 	output [PRO_ADDR_SPACE-1:0] pro_sram_waddr2, output [Q-1:0] pro_wbytemask2,
	output [Q*PRO_BW-1:0] pro_sram_wdata3, 	output [PRO_ADDR_SPACE-1:0] pro_sram_waddr3, output [Q-1:0] pro_wbytemask3,
	output [Q*PRO_BW-1:0] pro_sram_wdata4, 	output [PRO_ADDR_SPACE-1:0] pro_sram_waddr4, output [Q-1:0] pro_wbytemask4,
	output [Q*PRO_BW-1:0] pro_sram_wdata5, 	output [PRO_ADDR_SPACE-1:0] pro_sram_waddr5, output [Q-1:0] pro_wbytemask5,
	output [Q*PRO_BW-1:0] pro_sram_wdata6, 	output [PRO_ADDR_SPACE-1:0] pro_sram_waddr6, output [Q-1:0] pro_wbytemask6,
	output [Q*PRO_BW-1:0] pro_sram_wdata7, 	output [PRO_ADDR_SPACE-1:0] pro_sram_waddr7, output [Q-1:0] pro_wbytemask7,
	output [Q*PRO_BW-1:0] pro_sram_wdata8, 	output [PRO_ADDR_SPACE-1:0] pro_sram_waddr8, output [Q-1:0] pro_wbytemask8,
	output [Q*PRO_BW-1:0] pro_sram_wdata9, 	output [PRO_ADDR_SPACE-1:0] pro_sram_waddr9, output [Q-1:0] pro_wbytemask9,
	output [Q*PRO_BW-1:0] pro_sram_wdata10, output [PRO_ADDR_SPACE-1:0] pro_sram_waddr10, output [Q-1:0] pro_wbytemask10,
	output [Q*PRO_BW-1:0] pro_sram_wdata11, output [PRO_ADDR_SPACE-1:0] pro_sram_waddr11, output [Q-1:0] pro_wbytemask11,
	output [Q*PRO_BW-1:0] pro_sram_wdata12, output [PRO_ADDR_SPACE-1:0] pro_sram_waddr12, output [Q-1:0] pro_wbytemask12,
	output [Q*PRO_BW-1:0] pro_sram_wdata13, output [PRO_ADDR_SPACE-1:0] pro_sram_waddr13, output [Q-1:0] pro_wbytemask13,
	output [Q*PRO_BW-1:0] pro_sram_wdata14, output [PRO_ADDR_SPACE-1:0] pro_sram_waddr14, output [Q-1:0] pro_wbytemask14,
	output [Q*PRO_BW-1:0] pro_sram_wdata15, output [PRO_ADDR_SPACE-1:0] pro_sram_waddr15, output [Q-1:0] pro_wbytemask15,
	output reg part_finish
);

// ---- for master instance & declaration----
reg [3:0] iter, n_iter;
wire pingpong = iter[0]; // pingpong = 0 vid read from 0
wire [NEXT_ADDR_SPACE-1:0] next_sram_raddr_total; 
wire [VID_ADDR_SPACE-1:0] vid_sram_raddr_total;
assign next_sram_raddr0 = next_sram_raddr_total;	assign next_sram_raddr8 = next_sram_raddr_total;
assign next_sram_raddr1 = next_sram_raddr_total;	assign next_sram_raddr9 = next_sram_raddr_total;
assign next_sram_raddr2 = next_sram_raddr_total;	assign next_sram_raddr10 = next_sram_raddr_total;
assign next_sram_raddr3 = next_sram_raddr_total;	assign next_sram_raddr11 = next_sram_raddr_total;
assign next_sram_raddr4 = next_sram_raddr_total;	assign next_sram_raddr12 = next_sram_raddr_total;
assign next_sram_raddr5 = next_sram_raddr_total;	assign next_sram_raddr13 = next_sram_raddr_total;
assign next_sram_raddr6 = next_sram_raddr_total;	assign next_sram_raddr14 = next_sram_raddr_total;
assign next_sram_raddr7 = next_sram_raddr_total;	assign next_sram_raddr15 = next_sram_raddr_total;


assign pro_sram_raddr0 = next_sram_raddr_total; assign pro_sram_raddr8 = next_sram_raddr_total;
assign pro_sram_raddr1 = next_sram_raddr_total; assign pro_sram_raddr9 = next_sram_raddr_total;
assign pro_sram_raddr2 = next_sram_raddr_total; assign pro_sram_raddr10 = next_sram_raddr_total;
assign pro_sram_raddr3 = next_sram_raddr_total; assign pro_sram_raddr11 = next_sram_raddr_total;
assign pro_sram_raddr4 = next_sram_raddr_total; assign pro_sram_raddr12 = next_sram_raddr_total;
assign pro_sram_raddr5 = next_sram_raddr_total; assign pro_sram_raddr13 = next_sram_raddr_total;
assign pro_sram_raddr6 = next_sram_raddr_total; assign pro_sram_raddr14 = next_sram_raddr_total;
assign pro_sram_raddr7 = next_sram_raddr_total; assign pro_sram_raddr15 = next_sram_raddr_total;


// output 
wire master_finish;
wire [7:0] epoch, epoch_buff;
wire master_locsram_wen;
// input 
reg rst_n_master;
reg en_master;
// TODO mijs mjis 
reg [PRO_BW*K-1:0] in_mi_j; 
reg [PRO_BW*K-1:0] in_mj_i;
reg [7:0] batch_num, n_batch_num;
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr0;	wire [D*LOC_BW-1:0] master_loc_sram_wdata0;		wire [D-1:0] master_loc_wbytemask0;
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr1;	wire [D*LOC_BW-1:0] master_loc_sram_wdata1;		wire [D-1:0] master_loc_wbytemask1;
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr2;	wire [D*LOC_BW-1:0] master_loc_sram_wdata2;		wire [D-1:0] master_loc_wbytemask2;
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr3;	wire [D*LOC_BW-1:0] master_loc_sram_wdata3;		wire [D-1:0] master_loc_wbytemask3;
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr4;	wire [D*LOC_BW-1:0] master_loc_sram_wdata4;		wire [D-1:0] master_loc_wbytemask4;
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr5;	wire [D*LOC_BW-1:0] master_loc_sram_wdata5;		wire [D-1:0] master_loc_wbytemask5;
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr6;	wire [D*LOC_BW-1:0] master_loc_sram_wdata6;		wire [D-1:0] master_loc_wbytemask6;
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr7;	wire [D*LOC_BW-1:0] master_loc_sram_wdata7;		wire [D-1:0] master_loc_wbytemask7;
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr8;	wire [D*LOC_BW-1:0] master_loc_sram_wdata8;		wire [D-1:0] master_loc_wbytemask8;
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr9;	wire [D*LOC_BW-1:0] master_loc_sram_wdata9;		wire [D-1:0] master_loc_wbytemask9;
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr10;	wire [D*LOC_BW-1:0] master_loc_sram_wdata10;	wire [D-1:0] master_loc_wbytemask10;	
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr11;	wire [D*LOC_BW-1:0] master_loc_sram_wdata11;	wire [D-1:0] master_loc_wbytemask11;	
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr12;	wire [D*LOC_BW-1:0] master_loc_sram_wdata12;	wire [D-1:0] master_loc_wbytemask12;	
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr13;	wire [D*LOC_BW-1:0] master_loc_sram_wdata13;	wire [D-1:0] master_loc_wbytemask13;	
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr14;	wire [D*LOC_BW-1:0] master_loc_sram_wdata14;	wire [D-1:0] master_loc_wbytemask14;	
wire [LOC_ADDR_SPACE-1:0] master_loc_sram_waddr15;	wire [D*LOC_BW-1:0] master_loc_sram_wdata15;	wire [D-1:0] master_loc_wbytemask15;	
reg [3:0] tmpwaddr, n_tmpwaddr;
reg interfinish, n_interfinish;
parameter IDLE = 2'd0, WORKER = 2'd1, MASTER = 2'd2, FIN = 2'd3;
reg [1:0] state, n_state;

master_top_sram #(
.Q(Q),
.PRO_BW(PRO_BW),
.NEXT_BW(NEXT_BW),
.K(K),
.VID_BW(VID_BW),
.BUF_BW(5),
.OFFSET_BW(5),
.VID_ADDR_SPACE(VID_ADDR_SPACE),
.LOC_BW(LOC_BW),
.D(D),
.LOC_ADDR_SPACE(LOC_ADDR_SPACE),
.NEXT_ADDR_SPACE(NEXT_ADDR_SPACE),
.PRO_ADDR_SPACE(PRO_ADDR_SPACE)
) master_instn (
    .clk(clk),
    .enable_in(en_master),
    .rst_n_in(rst_n_master),
    .next_sram_rdata0(next_sram_rdata0), .next_sram_rdata8(next_sram_rdata8),
    .next_sram_rdata1(next_sram_rdata1), .next_sram_rdata9(next_sram_rdata9),
    .next_sram_rdata2(next_sram_rdata2), .next_sram_rdata10(next_sram_rdata10),
    .next_sram_rdata3(next_sram_rdata3), .next_sram_rdata11(next_sram_rdata11),
    .next_sram_rdata4(next_sram_rdata4), .next_sram_rdata12(next_sram_rdata12),
    .next_sram_rdata5(next_sram_rdata5), .next_sram_rdata13(next_sram_rdata13),
    .next_sram_rdata6(next_sram_rdata6), .next_sram_rdata14(next_sram_rdata14),
    .next_sram_rdata7(next_sram_rdata7), .next_sram_rdata15(next_sram_rdata15),
    
    .proposal_sram_rdata0(pro_sram_rdata0), .proposal_sram_rdata8(pro_sram_rdata8),
    .proposal_sram_rdata1(pro_sram_rdata1), .proposal_sram_rdata9(pro_sram_rdata9),
    .proposal_sram_rdata2(pro_sram_rdata2), .proposal_sram_rdata10(pro_sram_rdata10),
    .proposal_sram_rdata3(pro_sram_rdata3), .proposal_sram_rdata11(pro_sram_rdata11),
    .proposal_sram_rdata4(pro_sram_rdata4), .proposal_sram_rdata12(pro_sram_rdata12),
    .proposal_sram_rdata5(pro_sram_rdata5), .proposal_sram_rdata13(pro_sram_rdata13),
    .proposal_sram_rdata6(pro_sram_rdata6), .proposal_sram_rdata14(pro_sram_rdata14),
    .proposal_sram_rdata7(pro_sram_rdata7), .proposal_sram_rdata15(pro_sram_rdata15),
    
    .vid_sram_rdata0(vid_sram_rdata0),        .vid_sram_rdata8(vid_sram_rdata8),
    .vid_sram_rdata1(vid_sram_rdata1),        .vid_sram_rdata9(vid_sram_rdata9),
    .vid_sram_rdata2(vid_sram_rdata2),        .vid_sram_rdata10(vid_sram_rdata10),
    .vid_sram_rdata3(vid_sram_rdata3),        .vid_sram_rdata11(vid_sram_rdata11),
    .vid_sram_rdata4(vid_sram_rdata4),        .vid_sram_rdata12(vid_sram_rdata12),
    .vid_sram_rdata5(vid_sram_rdata5),        .vid_sram_rdata13(vid_sram_rdata13),
    .vid_sram_rdata6(vid_sram_rdata6),        .vid_sram_rdata14(vid_sram_rdata14),
    .vid_sram_rdata7(vid_sram_rdata7),        .vid_sram_rdata15(vid_sram_rdata15),

    .in_mi_j(in_mi_j),
    .in_mj_i(in_mj_i),
    .pingpong(pingpong),
    // output 
    .next_sram_raddr(next_sram_raddr_total), // same as proposal read addr
    .vid_sram_raddr(vid_sram_raddr_total),
    .epoch(epoch),
	.epoch_buff(epoch_buff),
    .vidsram_wen(vidsram_wen),
    .locsram_wen(master_locsram_wen), 
    .finish(master_finish),
    .vid_sram_wdata0(vid_sram_wdata0),     .vid_sram_waddr0(vid_sram_waddr0),
    .vid_sram_wdata1(vid_sram_wdata1),     .vid_sram_waddr1(vid_sram_waddr1),
    .vid_sram_wdata2(vid_sram_wdata2),     .vid_sram_waddr2(vid_sram_waddr2),
    .vid_sram_wdata3(vid_sram_wdata3),     .vid_sram_waddr3(vid_sram_waddr3),
    .vid_sram_wdata4(vid_sram_wdata4),     .vid_sram_waddr4(vid_sram_waddr4),
    .vid_sram_wdata5(vid_sram_wdata5),     .vid_sram_waddr5(vid_sram_waddr5),
    .vid_sram_wdata6(vid_sram_wdata6),     .vid_sram_waddr6(vid_sram_waddr6),
    .vid_sram_wdata7(vid_sram_wdata7),     .vid_sram_waddr7(vid_sram_waddr7),
    .vid_sram_wdata8(vid_sram_wdata8),     .vid_sram_waddr8(vid_sram_waddr8),
    .vid_sram_wdata9(vid_sram_wdata9),     .vid_sram_waddr9(vid_sram_waddr9),
    .vid_sram_wdata10(vid_sram_wdata10),   .vid_sram_waddr10(vid_sram_waddr10),    
    .vid_sram_wdata11(vid_sram_wdata11),   .vid_sram_waddr11(vid_sram_waddr11),    
    .vid_sram_wdata12(vid_sram_wdata12),   .vid_sram_waddr12(vid_sram_waddr12),    
    .vid_sram_wdata13(vid_sram_wdata13),   .vid_sram_waddr13(vid_sram_waddr13),    
    .vid_sram_wdata14(vid_sram_wdata14),   .vid_sram_waddr14(vid_sram_waddr14),    
    .vid_sram_wdata15(vid_sram_wdata15),   .vid_sram_waddr15(vid_sram_waddr15),

    .loc_sram_wdata0(master_loc_sram_wdata0)   ,  .loc_sram_waddr0(master_loc_sram_waddr0)    , .locsram_wbytemask0(master_loc_wbytemask0),
    .loc_sram_wdata1(master_loc_sram_wdata1)   ,  .loc_sram_waddr1(master_loc_sram_waddr1)    , .locsram_wbytemask1(master_loc_wbytemask1),
    .loc_sram_wdata2(master_loc_sram_wdata2)   ,  .loc_sram_waddr2(master_loc_sram_waddr2)    , .locsram_wbytemask2(master_loc_wbytemask2),
    .loc_sram_wdata3(master_loc_sram_wdata3)   ,  .loc_sram_waddr3(master_loc_sram_waddr3)    , .locsram_wbytemask3(master_loc_wbytemask3),
    .loc_sram_wdata4(master_loc_sram_wdata4)   ,  .loc_sram_waddr4(master_loc_sram_waddr4)    , .locsram_wbytemask4(master_loc_wbytemask4),
    .loc_sram_wdata5(master_loc_sram_wdata5)   ,  .loc_sram_waddr5(master_loc_sram_waddr5)    , .locsram_wbytemask5(master_loc_wbytemask5),
    .loc_sram_wdata6(master_loc_sram_wdata6)   ,  .loc_sram_waddr6(master_loc_sram_waddr6)    , .locsram_wbytemask6(master_loc_wbytemask6),
    .loc_sram_wdata7(master_loc_sram_wdata7)   ,  .loc_sram_waddr7(master_loc_sram_waddr7)    , .locsram_wbytemask7(master_loc_wbytemask7),
    .loc_sram_wdata8(master_loc_sram_wdata8)   ,  .loc_sram_waddr8(master_loc_sram_waddr8)    , .locsram_wbytemask8(master_loc_wbytemask8),
    .loc_sram_wdata9(master_loc_sram_wdata9)   ,  .loc_sram_waddr9(master_loc_sram_waddr9)    , .locsram_wbytemask9(master_loc_wbytemask9),
    .loc_sram_wdata10(master_loc_sram_wdata10) ,  .loc_sram_waddr10(master_loc_sram_waddr10)  , .locsram_wbytemask10(master_loc_wbytemask10),
    .loc_sram_wdata11(master_loc_sram_wdata11) ,  .loc_sram_waddr11(master_loc_sram_waddr11)  , .locsram_wbytemask11(master_loc_wbytemask11),
    .loc_sram_wdata12(master_loc_sram_wdata12) ,  .loc_sram_waddr12(master_loc_sram_waddr12)  , .locsram_wbytemask12(master_loc_wbytemask12),
    .loc_sram_wdata13(master_loc_sram_wdata13) ,  .loc_sram_waddr13(master_loc_sram_waddr13)  , .locsram_wbytemask13(master_loc_wbytemask13),
    .loc_sram_wdata14(master_loc_sram_wdata14) ,  .loc_sram_waddr14(master_loc_sram_waddr14)  , .locsram_wbytemask14(master_loc_wbytemask14),
    .loc_sram_wdata15(master_loc_sram_wdata15) ,  .loc_sram_waddr15(master_loc_sram_waddr15)  , .locsram_wbytemask15(master_loc_wbytemask15)
);
//---------------------------------------------

// all wires for worker_0~15 instances
reg en_worker, rst_n_worker;
wire [Q*VID_BW-1:0] w0_vid_rdata, w1_vid_rdata, w2_vid_rdata, w3_vid_rdata, w4_vid_rdata, w5_vid_rdata, w6_vid_rdata, w7_vid_rdata, w8_vid_rdata, w9_vid_rdata, w10_vid_rdata, w11_vid_rdata, w12_vid_rdata, w13_vid_rdata, w14_vid_rdata, w15_vid_rdata;
wire [D*DIST_BW-1:0] w0_dist_rdata, w1_dist_rdata, w2_dist_rdata, w3_dist_rdata, w4_dist_rdata, w5_dist_rdata, w6_dist_rdata, w7_dist_rdata, w8_dist_rdata, w9_dist_rdata, w10_dist_rdata, w11_dist_rdata, w12_dist_rdata, w13_dist_rdata, w14_dist_rdata, w15_dist_rdata;
wire [D*(LOC_BW-1)-1:0] w0_loc_rdata, w1_loc_rdata, w2_loc_rdata, w3_loc_rdata, w4_loc_rdata, w5_loc_rdata, w6_loc_rdata, w7_loc_rdata, w8_loc_rdata, w9_loc_rdata, w10_loc_rdata, w11_loc_rdata, w12_loc_rdata, w13_loc_rdata, w14_loc_rdata, w15_loc_rdata;

wire [3:0] sub_bat0, sub_bat1, sub_bat2, sub_bat3, sub_bat4, sub_bat5, sub_bat6, sub_bat7, sub_bat8, sub_bat9, sub_bat10, sub_bat11, sub_bat12, sub_bat13, sub_bat14, sub_bat15;
wire [VID_BW-1:0] vid0, vid1, vid2, vid3, vid4, vid5, vid6, vid7, vid8, vid9, vid10, vid11, vid12, vid13, vid14, vid15;
wire [Q-1:0] w0_next_bytemask, w1_next_bytemask, w2_next_bytemask, w3_next_bytemask, w4_next_bytemask, w5_next_bytemask, w6_next_bytemask, w7_next_bytemask, w8_next_bytemask, w9_next_bytemask, w10_next_bytemask, w11_next_bytemask, w12_next_bytemask, w13_next_bytemask, w14_next_bytemask, w15_next_bytemask;
wire [Q*NEXT_BW-1:0] w0_next_wdata, w1_next_wdata, w2_next_wdata, w3_next_wdata, w4_next_wdata, w5_next_wdata, w6_next_wdata, w7_next_wdata, w8_next_wdata, w9_next_wdata, w10_next_wdata, w11_next_wdata, w12_next_wdata, w13_next_wdata, w14_next_wdata, w15_next_wdata;
wire [NEXT_ADDR_SPACE-1:0] w0_next_waddr, w1_next_waddr, w2_next_waddr, w3_next_waddr, w4_next_waddr, w5_next_waddr, w6_next_waddr, w7_next_waddr, w8_next_waddr, w9_next_waddr, w10_next_waddr, w11_next_waddr, w12_next_waddr, w13_next_waddr, w14_next_waddr, w15_next_waddr;
wire [Q-1:0] w0_pro_bytemask, w1_pro_bytemask, w2_pro_bytemask, w3_pro_bytemask, w4_pro_bytemask, w5_pro_bytemask, w6_pro_bytemask, w7_pro_bytemask, w8_pro_bytemask, w9_pro_bytemask, w10_pro_bytemask, w11_pro_bytemask, w12_pro_bytemask, w13_pro_bytemask, w14_pro_bytemask, w15_pro_bytemask;
wire [Q*PRO_BW-1:0] w0_pro_wdata, w1_pro_wdata, w2_pro_wdata, w3_pro_wdata, w4_pro_wdata, w5_pro_wdata, w6_pro_wdata, w7_pro_wdata, w8_pro_wdata, w9_pro_wdata, w10_pro_wdata, w11_pro_wdata, w12_pro_wdata, w13_pro_wdata, w14_pro_wdata, w15_pro_wdata;
wire [PRO_ADDR_SPACE-1:0] w0_pro_waddr, w1_pro_waddr, w2_pro_waddr, w3_pro_waddr, w4_pro_waddr, w5_pro_waddr, w6_pro_waddr, w7_pro_waddr, w8_pro_waddr, w9_pro_waddr, w10_pro_waddr, w11_pro_waddr, w12_pro_waddr, w13_pro_waddr, w14_pro_waddr, w15_pro_waddr;
wire batch_finish0, batch_finish1, batch_finish2, batch_finish3, batch_finish4, batch_finish5, batch_finish6, batch_finish7, batch_finish8, batch_finish9, batch_finish10, batch_finish11, batch_finish12, batch_finish13, batch_finish14, batch_finish15;

wire [7:0] w0_proposal_num0, w0_proposal_num1, w0_proposal_num2, w0_proposal_num3, w0_proposal_num4, w0_proposal_num5, w0_proposal_num6, w0_proposal_num7, w0_proposal_num8, w0_proposal_num9, w0_proposal_num10, w0_proposal_num11, w0_proposal_num12, w0_proposal_num13, w0_proposal_num14, w0_proposal_num15;
wire [7:0] w1_proposal_num0, w1_proposal_num1, w1_proposal_num2, w1_proposal_num3, w1_proposal_num4, w1_proposal_num5, w1_proposal_num6, w1_proposal_num7, w1_proposal_num8, w1_proposal_num9, w1_proposal_num10, w1_proposal_num11, w1_proposal_num12, w1_proposal_num13, w1_proposal_num14, w1_proposal_num15;
wire [7:0] w2_proposal_num0, w2_proposal_num1, w2_proposal_num2, w2_proposal_num3, w2_proposal_num4, w2_proposal_num5, w2_proposal_num6, w2_proposal_num7, w2_proposal_num8, w2_proposal_num9, w2_proposal_num10, w2_proposal_num11, w2_proposal_num12, w2_proposal_num13, w2_proposal_num14, w2_proposal_num15;
wire [7:0] w3_proposal_num0, w3_proposal_num1, w3_proposal_num2, w3_proposal_num3, w3_proposal_num4, w3_proposal_num5, w3_proposal_num6, w3_proposal_num7, w3_proposal_num8, w3_proposal_num9, w3_proposal_num10, w3_proposal_num11, w3_proposal_num12, w3_proposal_num13, w3_proposal_num14, w3_proposal_num15;
wire [7:0] w4_proposal_num0, w4_proposal_num1, w4_proposal_num2, w4_proposal_num3, w4_proposal_num4, w4_proposal_num5, w4_proposal_num6, w4_proposal_num7, w4_proposal_num8, w4_proposal_num9, w4_proposal_num10, w4_proposal_num11, w4_proposal_num12, w4_proposal_num13, w4_proposal_num14, w4_proposal_num15;
wire [7:0] w5_proposal_num0, w5_proposal_num1, w5_proposal_num2, w5_proposal_num3, w5_proposal_num4, w5_proposal_num5, w5_proposal_num6, w5_proposal_num7, w5_proposal_num8, w5_proposal_num9, w5_proposal_num10, w5_proposal_num11, w5_proposal_num12, w5_proposal_num13, w5_proposal_num14, w5_proposal_num15;
wire [7:0] w6_proposal_num0, w6_proposal_num1, w6_proposal_num2, w6_proposal_num3, w6_proposal_num4, w6_proposal_num5, w6_proposal_num6, w6_proposal_num7, w6_proposal_num8, w6_proposal_num9, w6_proposal_num10, w6_proposal_num11, w6_proposal_num12, w6_proposal_num13, w6_proposal_num14, w6_proposal_num15;
wire [7:0] w7_proposal_num0, w7_proposal_num1, w7_proposal_num2, w7_proposal_num3, w7_proposal_num4, w7_proposal_num5, w7_proposal_num6, w7_proposal_num7, w7_proposal_num8, w7_proposal_num9, w7_proposal_num10, w7_proposal_num11, w7_proposal_num12, w7_proposal_num13, w7_proposal_num14, w7_proposal_num15;
wire [7:0] w8_proposal_num0, w8_proposal_num1, w8_proposal_num2, w8_proposal_num3, w8_proposal_num4, w8_proposal_num5, w8_proposal_num6, w8_proposal_num7, w8_proposal_num8, w8_proposal_num9, w8_proposal_num10, w8_proposal_num11, w8_proposal_num12, w8_proposal_num13, w8_proposal_num14, w8_proposal_num15;
wire [7:0] w9_proposal_num0, w9_proposal_num1, w9_proposal_num2, w9_proposal_num3, w9_proposal_num4, w9_proposal_num5, w9_proposal_num6, w9_proposal_num7, w9_proposal_num8, w9_proposal_num9, w9_proposal_num10, w9_proposal_num11, w9_proposal_num12, w9_proposal_num13, w9_proposal_num14, w9_proposal_num15;
wire [7:0] w10_proposal_num0, w10_proposal_num1, w10_proposal_num2, w10_proposal_num3, w10_proposal_num4, w10_proposal_num5, w10_proposal_num6, w10_proposal_num7, w10_proposal_num8, w10_proposal_num9, w10_proposal_num10, w10_proposal_num11, w10_proposal_num12, w10_proposal_num13, w10_proposal_num14, w10_proposal_num15;
wire [7:0] w11_proposal_num0, w11_proposal_num1, w11_proposal_num2, w11_proposal_num3, w11_proposal_num4, w11_proposal_num5, w11_proposal_num6, w11_proposal_num7, w11_proposal_num8, w11_proposal_num9, w11_proposal_num10, w11_proposal_num11, w11_proposal_num12, w11_proposal_num13, w11_proposal_num14, w11_proposal_num15;
wire [7:0] w12_proposal_num0, w12_proposal_num1, w12_proposal_num2, w12_proposal_num3, w12_proposal_num4, w12_proposal_num5, w12_proposal_num6, w12_proposal_num7, w12_proposal_num8, w12_proposal_num9, w12_proposal_num10, w12_proposal_num11, w12_proposal_num12, w12_proposal_num13, w12_proposal_num14, w12_proposal_num15;
wire [7:0] w13_proposal_num0, w13_proposal_num1, w13_proposal_num2, w13_proposal_num3, w13_proposal_num4, w13_proposal_num5, w13_proposal_num6, w13_proposal_num7, w13_proposal_num8, w13_proposal_num9, w13_proposal_num10, w13_proposal_num11, w13_proposal_num12, w13_proposal_num13, w13_proposal_num14, w13_proposal_num15;
wire [7:0] w14_proposal_num0, w14_proposal_num1, w14_proposal_num2, w14_proposal_num3, w14_proposal_num4, w14_proposal_num5, w14_proposal_num6, w14_proposal_num7, w14_proposal_num8, w14_proposal_num9, w14_proposal_num10, w14_proposal_num11, w14_proposal_num12, w14_proposal_num13, w14_proposal_num14, w14_proposal_num15;
wire [7:0] w15_proposal_num0, w15_proposal_num1, w15_proposal_num2, w15_proposal_num3, w15_proposal_num4, w15_proposal_num5, w15_proposal_num6, w15_proposal_num7, w15_proposal_num8, w15_proposal_num9, w15_proposal_num10, w15_proposal_num11, w15_proposal_num12, w15_proposal_num13, w15_proposal_num14, w15_proposal_num15;


worker #(.WORK_IDX(0)) worker_0
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w0_vid_rdata),
	.dist_rdata(w0_dist_rdata),
	.loc_rdata(w0_loc_rdata),

	.sub_bat(sub_bat0),
	.vid(vid0),
	.next_bytemask(w0_next_bytemask),
	.next_wdata(w0_next_wdata),
	.next_waddr(w0_next_waddr),
	.pro_bytemask(w0_pro_bytemask),
	.pro_wdata(w0_pro_wdata),
	.pro_waddr(w0_pro_waddr),
	.ready(),
	.batch_finish(batch_finish0),
	.wen_delay(wen0),
	.proposal_num0(w0_proposal_num0),
	.proposal_num1(w0_proposal_num1),
	.proposal_num2(w0_proposal_num2),
	.proposal_num3(w0_proposal_num3),
	.proposal_num4(w0_proposal_num4),
	.proposal_num5(w0_proposal_num5),
	.proposal_num6(w0_proposal_num6),
	.proposal_num7(w0_proposal_num7),
	.proposal_num8(w0_proposal_num8),
	.proposal_num9(w0_proposal_num9),
	.proposal_num10(w0_proposal_num10),
	.proposal_num11(w0_proposal_num11),
	.proposal_num12(w0_proposal_num12),
	.proposal_num13(w0_proposal_num13),
	.proposal_num14(w0_proposal_num14),
	.proposal_num15(w0_proposal_num15)
);

worker #(.WORK_IDX(1)) worker_1
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w1_vid_rdata),
	.dist_rdata(w1_dist_rdata),
	.loc_rdata(w1_loc_rdata),

	.sub_bat(sub_bat1),
	.vid(vid1),
	.next_bytemask(w1_next_bytemask),
	.next_wdata(w1_next_wdata),
	.next_waddr(w1_next_waddr),
	.pro_bytemask(w1_pro_bytemask),
	.pro_wdata(w1_pro_wdata),
	.pro_waddr(w1_pro_waddr),
	.ready(),
	.batch_finish(batch_finish1),
	.wen_delay(wen1),
	.proposal_num0(w1_proposal_num0),
	.proposal_num1(w1_proposal_num1),
	.proposal_num2(w1_proposal_num2),
	.proposal_num3(w1_proposal_num3),
	.proposal_num4(w1_proposal_num4),
	.proposal_num5(w1_proposal_num5),
	.proposal_num6(w1_proposal_num6),
	.proposal_num7(w1_proposal_num7),
	.proposal_num8(w1_proposal_num8),
	.proposal_num9(w1_proposal_num9),
	.proposal_num10(w1_proposal_num10),
	.proposal_num11(w1_proposal_num11),
	.proposal_num12(w1_proposal_num12),
	.proposal_num13(w1_proposal_num13),
	.proposal_num14(w1_proposal_num14),
	.proposal_num15(w1_proposal_num15)
);

worker #(.WORK_IDX(2)) worker_2
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w2_vid_rdata),
	.dist_rdata(w2_dist_rdata),
	.loc_rdata(w2_loc_rdata),

	.sub_bat(sub_bat2),
	.vid(vid2),
	.next_bytemask(w2_next_bytemask),
	.next_wdata(w2_next_wdata),
	.next_waddr(w2_next_waddr),
	.pro_bytemask(w2_pro_bytemask),
	.pro_wdata(w2_pro_wdata),
	.pro_waddr(w2_pro_waddr),
	.ready(),
	.batch_finish(batch_finish2),
	.wen_delay(wen2),
	.proposal_num0(w2_proposal_num0),
	.proposal_num1(w2_proposal_num1),
	.proposal_num2(w2_proposal_num2),
	.proposal_num3(w2_proposal_num3),
	.proposal_num4(w2_proposal_num4),
	.proposal_num5(w2_proposal_num5),
	.proposal_num6(w2_proposal_num6),
	.proposal_num7(w2_proposal_num7),
	.proposal_num8(w2_proposal_num8),
	.proposal_num9(w2_proposal_num9),
	.proposal_num10(w2_proposal_num10),
	.proposal_num11(w2_proposal_num11),
	.proposal_num12(w2_proposal_num12),
	.proposal_num13(w2_proposal_num13),
	.proposal_num14(w2_proposal_num14),
	.proposal_num15(w2_proposal_num15)
);

worker #(.WORK_IDX(3)) worker_3
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w3_vid_rdata),
	.dist_rdata(w3_dist_rdata),
	.loc_rdata(w3_loc_rdata),

	.sub_bat(sub_bat3),
	.vid(vid3),
	.next_bytemask(w3_next_bytemask),
	.next_wdata(w3_next_wdata),
	.next_waddr(w3_next_waddr),
	.pro_bytemask(w3_pro_bytemask),
	.pro_wdata(w3_pro_wdata),
	.pro_waddr(w3_pro_waddr),
	.ready(),
	.batch_finish(batch_finish3),
	.wen_delay(wen3),
	.proposal_num0(w3_proposal_num0),
	.proposal_num1(w3_proposal_num1),
	.proposal_num2(w3_proposal_num2),
	.proposal_num3(w3_proposal_num3),
	.proposal_num4(w3_proposal_num4),
	.proposal_num5(w3_proposal_num5),
	.proposal_num6(w3_proposal_num6),
	.proposal_num7(w3_proposal_num7),
	.proposal_num8(w3_proposal_num8),
	.proposal_num9(w3_proposal_num9),
	.proposal_num10(w3_proposal_num10),
	.proposal_num11(w3_proposal_num11),
	.proposal_num12(w3_proposal_num12),
	.proposal_num13(w3_proposal_num13),
	.proposal_num14(w3_proposal_num14),
	.proposal_num15(w3_proposal_num15)
);

worker #(.WORK_IDX(4)) worker_4
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w4_vid_rdata),
	.dist_rdata(w4_dist_rdata),
	.loc_rdata(w4_loc_rdata),

	.sub_bat(sub_bat4),
	.vid(vid4),
	.next_bytemask(w4_next_bytemask),
	.next_wdata(w4_next_wdata),
	.next_waddr(w4_next_waddr),
	.pro_bytemask(w4_pro_bytemask),
	.pro_wdata(w4_pro_wdata),
	.pro_waddr(w4_pro_waddr),
	.ready(),
	.batch_finish(batch_finish4),
	.wen_delay(wen4),
	.proposal_num0(w4_proposal_num0),
	.proposal_num1(w4_proposal_num1),
	.proposal_num2(w4_proposal_num2),
	.proposal_num3(w4_proposal_num3),
	.proposal_num4(w4_proposal_num4),
	.proposal_num5(w4_proposal_num5),
	.proposal_num6(w4_proposal_num6),
	.proposal_num7(w4_proposal_num7),
	.proposal_num8(w4_proposal_num8),
	.proposal_num9(w4_proposal_num9),
	.proposal_num10(w4_proposal_num10),
	.proposal_num11(w4_proposal_num11),
	.proposal_num12(w4_proposal_num12),
	.proposal_num13(w4_proposal_num13),
	.proposal_num14(w4_proposal_num14),
	.proposal_num15(w4_proposal_num15)
);

worker #(.WORK_IDX(5)) worker_5
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w5_vid_rdata),
	.dist_rdata(w5_dist_rdata),
	.loc_rdata(w5_loc_rdata),

	.sub_bat(sub_bat5),
	.vid(vid5),
	.next_bytemask(w5_next_bytemask),
	.next_wdata(w5_next_wdata),
	.next_waddr(w5_next_waddr),
	.pro_bytemask(w5_pro_bytemask),
	.pro_wdata(w5_pro_wdata),
	.pro_waddr(w5_pro_waddr),
	.ready(),
	.batch_finish(batch_finish5),
	.wen_delay(wen5),
	.proposal_num0(w5_proposal_num0),
	.proposal_num1(w5_proposal_num1),
	.proposal_num2(w5_proposal_num2),
	.proposal_num3(w5_proposal_num3),
	.proposal_num4(w5_proposal_num4),
	.proposal_num5(w5_proposal_num5),
	.proposal_num6(w5_proposal_num6),
	.proposal_num7(w5_proposal_num7),
	.proposal_num8(w5_proposal_num8),
	.proposal_num9(w5_proposal_num9),
	.proposal_num10(w5_proposal_num10),
	.proposal_num11(w5_proposal_num11),
	.proposal_num12(w5_proposal_num12),
	.proposal_num13(w5_proposal_num13),
	.proposal_num14(w5_proposal_num14),
	.proposal_num15(w5_proposal_num15)
);

worker #(.WORK_IDX(6)) worker_6
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w6_vid_rdata),
	.dist_rdata(w6_dist_rdata),
	.loc_rdata(w6_loc_rdata),

	.sub_bat(sub_bat6),
	.vid(vid6),
	.next_bytemask(w6_next_bytemask),
	.next_wdata(w6_next_wdata),
	.next_waddr(w6_next_waddr),
	.pro_bytemask(w6_pro_bytemask),
	.pro_wdata(w6_pro_wdata),
	.pro_waddr(w6_pro_waddr),
	.ready(),
	.batch_finish(batch_finish6),
	.wen_delay(wen6),
	.proposal_num0(w6_proposal_num0),
	.proposal_num1(w6_proposal_num1),
	.proposal_num2(w6_proposal_num2),
	.proposal_num3(w6_proposal_num3),
	.proposal_num4(w6_proposal_num4),
	.proposal_num5(w6_proposal_num5),
	.proposal_num6(w6_proposal_num6),
	.proposal_num7(w6_proposal_num7),
	.proposal_num8(w6_proposal_num8),
	.proposal_num9(w6_proposal_num9),
	.proposal_num10(w6_proposal_num10),
	.proposal_num11(w6_proposal_num11),
	.proposal_num12(w6_proposal_num12),
	.proposal_num13(w6_proposal_num13),
	.proposal_num14(w6_proposal_num14),
	.proposal_num15(w6_proposal_num15)
);

worker #(.WORK_IDX(7)) worker_7
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w7_vid_rdata),
	.dist_rdata(w7_dist_rdata),
	.loc_rdata(w7_loc_rdata),

	.sub_bat(sub_bat7),
	.vid(vid7),
	.next_bytemask(w7_next_bytemask),
	.next_wdata(w7_next_wdata),
	.next_waddr(w7_next_waddr),
	.pro_bytemask(w7_pro_bytemask),
	.pro_wdata(w7_pro_wdata),
	.pro_waddr(w7_pro_waddr),
	.ready(),
	.batch_finish(batch_finish7),
	.wen_delay(wen7),
	.proposal_num0(w7_proposal_num0),
	.proposal_num1(w7_proposal_num1),
	.proposal_num2(w7_proposal_num2),
	.proposal_num3(w7_proposal_num3),
	.proposal_num4(w7_proposal_num4),
	.proposal_num5(w7_proposal_num5),
	.proposal_num6(w7_proposal_num6),
	.proposal_num7(w7_proposal_num7),
	.proposal_num8(w7_proposal_num8),
	.proposal_num9(w7_proposal_num9),
	.proposal_num10(w7_proposal_num10),
	.proposal_num11(w7_proposal_num11),
	.proposal_num12(w7_proposal_num12),
	.proposal_num13(w7_proposal_num13),
	.proposal_num14(w7_proposal_num14),
	.proposal_num15(w7_proposal_num15)
);

worker #(.WORK_IDX(8)) worker_8
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w8_vid_rdata),
	.dist_rdata(w8_dist_rdata),
	.loc_rdata(w8_loc_rdata),

	.sub_bat(sub_bat8),
	.vid(vid8),
	.next_bytemask(w8_next_bytemask),
	.next_wdata(w8_next_wdata),
	.next_waddr(w8_next_waddr),
	.pro_bytemask(w8_pro_bytemask),
	.pro_wdata(w8_pro_wdata),
	.pro_waddr(w8_pro_waddr),
	.ready(),
	.batch_finish(batch_finish8),
	.wen_delay(wen8),
	.proposal_num0(w8_proposal_num0),
	.proposal_num1(w8_proposal_num1),
	.proposal_num2(w8_proposal_num2),
	.proposal_num3(w8_proposal_num3),
	.proposal_num4(w8_proposal_num4),
	.proposal_num5(w8_proposal_num5),
	.proposal_num6(w8_proposal_num6),
	.proposal_num7(w8_proposal_num7),
	.proposal_num8(w8_proposal_num8),
	.proposal_num9(w8_proposal_num9),
	.proposal_num10(w8_proposal_num10),
	.proposal_num11(w8_proposal_num11),
	.proposal_num12(w8_proposal_num12),
	.proposal_num13(w8_proposal_num13),
	.proposal_num14(w8_proposal_num14),
	.proposal_num15(w8_proposal_num15)
);

worker #(.WORK_IDX(9)) worker_9
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w9_vid_rdata),
	.dist_rdata(w9_dist_rdata),
	.loc_rdata(w9_loc_rdata),

	.sub_bat(sub_bat9),
	.vid(vid9),
	.next_bytemask(w9_next_bytemask),
	.next_wdata(w9_next_wdata),
	.next_waddr(w9_next_waddr),
	.pro_bytemask(w9_pro_bytemask),
	.pro_wdata(w9_pro_wdata),
	.pro_waddr(w9_pro_waddr),
	.ready(),
	.batch_finish(batch_finish9),
	.wen_delay(wen9),
	.proposal_num0(w9_proposal_num0),
	.proposal_num1(w9_proposal_num1),
	.proposal_num2(w9_proposal_num2),
	.proposal_num3(w9_proposal_num3),
	.proposal_num4(w9_proposal_num4),
	.proposal_num5(w9_proposal_num5),
	.proposal_num6(w9_proposal_num6),
	.proposal_num7(w9_proposal_num7),
	.proposal_num8(w9_proposal_num8),
	.proposal_num9(w9_proposal_num9),
	.proposal_num10(w9_proposal_num10),
	.proposal_num11(w9_proposal_num11),
	.proposal_num12(w9_proposal_num12),
	.proposal_num13(w9_proposal_num13),
	.proposal_num14(w9_proposal_num14),
	.proposal_num15(w9_proposal_num15)
);

worker #(.WORK_IDX(10)) worker_10
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w10_vid_rdata),
	.dist_rdata(w10_dist_rdata),
	.loc_rdata(w10_loc_rdata),

	.sub_bat(sub_bat10),
	.vid(vid10),
	.next_bytemask(w10_next_bytemask),
	.next_wdata(w10_next_wdata),
	.next_waddr(w10_next_waddr),
	.pro_bytemask(w10_pro_bytemask),
	.pro_wdata(w10_pro_wdata),
	.pro_waddr(w10_pro_waddr),
	.ready(),
	.batch_finish(batch_finish10),
	.wen_delay(wen10),
	.proposal_num0(w10_proposal_num0),
	.proposal_num1(w10_proposal_num1),
	.proposal_num2(w10_proposal_num2),
	.proposal_num3(w10_proposal_num3),
	.proposal_num4(w10_proposal_num4),
	.proposal_num5(w10_proposal_num5),
	.proposal_num6(w10_proposal_num6),
	.proposal_num7(w10_proposal_num7),
	.proposal_num8(w10_proposal_num8),
	.proposal_num9(w10_proposal_num9),
	.proposal_num10(w10_proposal_num10),
	.proposal_num11(w10_proposal_num11),
	.proposal_num12(w10_proposal_num12),
	.proposal_num13(w10_proposal_num13),
	.proposal_num14(w10_proposal_num14),
	.proposal_num15(w10_proposal_num15)
);

worker #(.WORK_IDX(11)) worker_11
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w11_vid_rdata),
	.dist_rdata(w11_dist_rdata),
	.loc_rdata(w11_loc_rdata),

	.sub_bat(sub_bat11),
	.vid(vid11),
	.next_bytemask(w11_next_bytemask),
	.next_wdata(w11_next_wdata),
	.next_waddr(w11_next_waddr),
	.pro_bytemask(w11_pro_bytemask),
	.pro_wdata(w11_pro_wdata),
	.pro_waddr(w11_pro_waddr),
	.ready(),
	.batch_finish(batch_finish11),
	.wen_delay(wen11),
	.proposal_num0(w11_proposal_num0),
	.proposal_num1(w11_proposal_num1),
	.proposal_num2(w11_proposal_num2),
	.proposal_num3(w11_proposal_num3),
	.proposal_num4(w11_proposal_num4),
	.proposal_num5(w11_proposal_num5),
	.proposal_num6(w11_proposal_num6),
	.proposal_num7(w11_proposal_num7),
	.proposal_num8(w11_proposal_num8),
	.proposal_num9(w11_proposal_num9),
	.proposal_num10(w11_proposal_num10),
	.proposal_num11(w11_proposal_num11),
	.proposal_num12(w11_proposal_num12),
	.proposal_num13(w11_proposal_num13),
	.proposal_num14(w11_proposal_num14),
	.proposal_num15(w11_proposal_num15)
);

worker #(.WORK_IDX(12)) worker_12
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w12_vid_rdata),
	.dist_rdata(w12_dist_rdata),
	.loc_rdata(w12_loc_rdata),

	.sub_bat(sub_bat12),
	.vid(vid12),
	.next_bytemask(w12_next_bytemask),
	.next_wdata(w12_next_wdata),
	.next_waddr(w12_next_waddr),
	.pro_bytemask(w12_pro_bytemask),
	.pro_wdata(w12_pro_wdata),
	.pro_waddr(w12_pro_waddr),
	.ready(),
	.batch_finish(batch_finish12),
	.wen_delay(wen12),
	.proposal_num0(w12_proposal_num0),
	.proposal_num1(w12_proposal_num1),
	.proposal_num2(w12_proposal_num2),
	.proposal_num3(w12_proposal_num3),
	.proposal_num4(w12_proposal_num4),
	.proposal_num5(w12_proposal_num5),
	.proposal_num6(w12_proposal_num6),
	.proposal_num7(w12_proposal_num7),
	.proposal_num8(w12_proposal_num8),
	.proposal_num9(w12_proposal_num9),
	.proposal_num10(w12_proposal_num10),
	.proposal_num11(w12_proposal_num11),
	.proposal_num12(w12_proposal_num12),
	.proposal_num13(w12_proposal_num13),
	.proposal_num14(w12_proposal_num14),
	.proposal_num15(w12_proposal_num15)
);

worker #(.WORK_IDX(13)) worker_13
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w13_vid_rdata),
	.dist_rdata(w13_dist_rdata),
	.loc_rdata(w13_loc_rdata),

	.sub_bat(sub_bat13),
	.vid(vid13),
	.next_bytemask(w13_next_bytemask),
	.next_wdata(w13_next_wdata),
	.next_waddr(w13_next_waddr),
	.pro_bytemask(w13_pro_bytemask),
	.pro_wdata(w13_pro_wdata),
	.pro_waddr(w13_pro_waddr),
	.ready(),
	.batch_finish(batch_finish13),
	.wen_delay(wen13),
	.proposal_num0(w13_proposal_num0),
	.proposal_num1(w13_proposal_num1),
	.proposal_num2(w13_proposal_num2),
	.proposal_num3(w13_proposal_num3),
	.proposal_num4(w13_proposal_num4),
	.proposal_num5(w13_proposal_num5),
	.proposal_num6(w13_proposal_num6),
	.proposal_num7(w13_proposal_num7),
	.proposal_num8(w13_proposal_num8),
	.proposal_num9(w13_proposal_num9),
	.proposal_num10(w13_proposal_num10),
	.proposal_num11(w13_proposal_num11),
	.proposal_num12(w13_proposal_num12),
	.proposal_num13(w13_proposal_num13),
	.proposal_num14(w13_proposal_num14),
	.proposal_num15(w13_proposal_num15)
);

worker #(.WORK_IDX(14)) worker_14
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w14_vid_rdata),
	.dist_rdata(w14_dist_rdata),
	.loc_rdata(w14_loc_rdata),

	.sub_bat(sub_bat14),
	.vid(vid14),
	.next_bytemask(w14_next_bytemask),
	.next_wdata(w14_next_wdata),
	.next_waddr(w14_next_waddr),
	.pro_bytemask(w14_pro_bytemask),
	.pro_wdata(w14_pro_wdata),
	.pro_waddr(w14_pro_waddr),
	.ready(),
	.batch_finish(batch_finish14),
	.wen_delay(wen14),
	.proposal_num0(w14_proposal_num0),
	.proposal_num1(w14_proposal_num1),
	.proposal_num2(w14_proposal_num2),
	.proposal_num3(w14_proposal_num3),
	.proposal_num4(w14_proposal_num4),
	.proposal_num5(w14_proposal_num5),
	.proposal_num6(w14_proposal_num6),
	.proposal_num7(w14_proposal_num7),
	.proposal_num8(w14_proposal_num8),
	.proposal_num9(w14_proposal_num9),
	.proposal_num10(w14_proposal_num10),
	.proposal_num11(w14_proposal_num11),
	.proposal_num12(w14_proposal_num12),
	.proposal_num13(w14_proposal_num13),
	.proposal_num14(w14_proposal_num14),
	.proposal_num15(w14_proposal_num15)
);

worker #(.WORK_IDX(15)) worker_15
(
	.clk(clk),
	.en(en_worker),
	.rst_n(rst_n_worker),
	.batch_num(batch_num),
	.vid_rdata(w15_vid_rdata),
	.dist_rdata(w15_dist_rdata),
	.loc_rdata(w15_loc_rdata),

	.sub_bat(sub_bat15),
	.vid(vid15),
	.next_bytemask(w15_next_bytemask),
	.next_wdata(w15_next_wdata),
	.next_waddr(w15_next_waddr),
	.pro_bytemask(w15_pro_bytemask),
	.pro_wdata(w15_pro_wdata),
	.pro_waddr(w15_pro_waddr),
	.ready(),
	.batch_finish(batch_finish15),
	.wen_delay(wen15),
	.proposal_num0(w15_proposal_num0),
	.proposal_num1(w15_proposal_num1),
	.proposal_num2(w15_proposal_num2),
	.proposal_num3(w15_proposal_num3),
	.proposal_num4(w15_proposal_num4),
	.proposal_num5(w15_proposal_num5),
	.proposal_num6(w15_proposal_num6),
	.proposal_num7(w15_proposal_num7),
	.proposal_num8(w15_proposal_num8),
	.proposal_num9(w15_proposal_num9),
	.proposal_num10(w15_proposal_num10),
	.proposal_num11(w15_proposal_num11),
	.proposal_num12(w15_proposal_num12),
	.proposal_num13(w15_proposal_num13),
	.proposal_num14(w15_proposal_num14),
	.proposal_num15(w15_proposal_num15)
);

assign worker_wen = (state == MASTER) ? 1'b0 : wen0;

// next_sram write out
assign next_wbytemask0 = w0_next_bytemask;
assign next_wbytemask1 = w1_next_bytemask;
assign next_wbytemask2 = w2_next_bytemask;
assign next_wbytemask3 = w3_next_bytemask;
assign next_wbytemask4 = w4_next_bytemask;
assign next_wbytemask5 = w5_next_bytemask;
assign next_wbytemask6 = w6_next_bytemask;
assign next_wbytemask7 = w7_next_bytemask;
assign next_wbytemask8 = w8_next_bytemask;
assign next_wbytemask9 = w9_next_bytemask;
assign next_wbytemask10 = w10_next_bytemask;
assign next_wbytemask11 = w11_next_bytemask;
assign next_wbytemask12 = w12_next_bytemask;
assign next_wbytemask13 = w13_next_bytemask;
assign next_wbytemask14 = w14_next_bytemask;
assign next_wbytemask15 = w15_next_bytemask;

assign next_sram_wdata0 = w0_next_wdata;
assign next_sram_wdata1 = w1_next_wdata;
assign next_sram_wdata2 = w2_next_wdata;
assign next_sram_wdata3 = w3_next_wdata;
assign next_sram_wdata4 = w4_next_wdata;
assign next_sram_wdata5 = w5_next_wdata;
assign next_sram_wdata6 = w6_next_wdata;
assign next_sram_wdata7 = w7_next_wdata;
assign next_sram_wdata8 = w8_next_wdata;
assign next_sram_wdata9 = w9_next_wdata;
assign next_sram_wdata10 = w10_next_wdata;
assign next_sram_wdata11 = w11_next_wdata;
assign next_sram_wdata12 = w12_next_wdata;
assign next_sram_wdata13 = w13_next_wdata;
assign next_sram_wdata14 = w14_next_wdata;
assign next_sram_wdata15 = w15_next_wdata;

assign next_sram_waddr0 = w0_next_waddr;
assign next_sram_waddr1 = w1_next_waddr;
assign next_sram_waddr2 = w2_next_waddr;
assign next_sram_waddr3 = w3_next_waddr;
assign next_sram_waddr4 = w4_next_waddr;
assign next_sram_waddr5 = w5_next_waddr;
assign next_sram_waddr6 = w6_next_waddr;
assign next_sram_waddr7 = w7_next_waddr;
assign next_sram_waddr8 = w8_next_waddr;
assign next_sram_waddr9 = w9_next_waddr;
assign next_sram_waddr10 = w10_next_waddr;
assign next_sram_waddr11 = w11_next_waddr;
assign next_sram_waddr12 = w12_next_waddr;
assign next_sram_waddr13 = w13_next_waddr;
assign next_sram_waddr14 = w14_next_waddr;
assign next_sram_waddr15 = w15_next_waddr;

// pro sram write out
assign pro_wbytemask0 = w0_pro_bytemask;
assign pro_wbytemask1 = w1_pro_bytemask;
assign pro_wbytemask2 = w2_pro_bytemask;
assign pro_wbytemask3 = w3_pro_bytemask;
assign pro_wbytemask4 = w4_pro_bytemask;
assign pro_wbytemask5 = w5_pro_bytemask;
assign pro_wbytemask6 = w6_pro_bytemask;
assign pro_wbytemask7 = w7_pro_bytemask;
assign pro_wbytemask8 = w8_pro_bytemask;
assign pro_wbytemask9 = w9_pro_bytemask;
assign pro_wbytemask10 = w10_pro_bytemask;
assign pro_wbytemask11 = w11_pro_bytemask;
assign pro_wbytemask12 = w12_pro_bytemask;
assign pro_wbytemask13 = w13_pro_bytemask;
assign pro_wbytemask14 = w14_pro_bytemask;
assign pro_wbytemask15 = w15_pro_bytemask;

assign pro_sram_wdata0 = w0_pro_wdata;
assign pro_sram_wdata1 = w1_pro_wdata;
assign pro_sram_wdata2 = w2_pro_wdata;
assign pro_sram_wdata3 = w3_pro_wdata;
assign pro_sram_wdata4 = w4_pro_wdata;
assign pro_sram_wdata5 = w5_pro_wdata;
assign pro_sram_wdata6 = w6_pro_wdata;
assign pro_sram_wdata7 = w7_pro_wdata;
assign pro_sram_wdata8 = w8_pro_wdata;
assign pro_sram_wdata9 = w9_pro_wdata;
assign pro_sram_wdata10 = w10_pro_wdata;
assign pro_sram_wdata11 = w11_pro_wdata;
assign pro_sram_wdata12 = w12_pro_wdata;
assign pro_sram_wdata13 = w13_pro_wdata;
assign pro_sram_wdata14 = w14_pro_wdata;
assign pro_sram_wdata15 = w15_pro_wdata;

assign pro_sram_waddr0 = w0_pro_waddr;
assign pro_sram_waddr1 = w1_pro_waddr;
assign pro_sram_waddr2 = w2_pro_waddr;
assign pro_sram_waddr3 = w3_pro_waddr;
assign pro_sram_waddr4 = w4_pro_waddr;
assign pro_sram_waddr5 = w5_pro_waddr;
assign pro_sram_waddr6 = w6_pro_waddr;
assign pro_sram_waddr7 = w7_pro_waddr;
assign pro_sram_waddr8 = w8_pro_waddr;
assign pro_sram_waddr9 = w9_pro_waddr;
assign pro_sram_waddr10 = w10_pro_waddr;
assign pro_sram_waddr11 = w11_pro_waddr;
assign pro_sram_waddr12 = w12_pro_waddr;
assign pro_sram_waddr13 = w13_pro_waddr;
assign pro_sram_waddr14 = w14_pro_waddr;
assign pro_sram_waddr15 = w15_pro_waddr;

// loc sram read in
assign loc_sram_raddr0 = sub_bat0;
assign loc_sram_raddr1 = sub_bat1;
assign loc_sram_raddr2 = sub_bat2;
assign loc_sram_raddr3 = sub_bat3;
assign loc_sram_raddr4 = sub_bat4;
assign loc_sram_raddr5 = sub_bat5;
assign loc_sram_raddr6 = sub_bat6;
assign loc_sram_raddr7 = sub_bat7;
assign loc_sram_raddr8 = sub_bat8;
assign loc_sram_raddr9 = sub_bat9;
assign loc_sram_raddr10 = sub_bat10;
assign loc_sram_raddr11 = sub_bat11;
assign loc_sram_raddr12 = sub_bat12;
assign loc_sram_raddr13 = sub_bat13;
assign loc_sram_raddr14 = sub_bat14;
assign loc_sram_raddr15 = sub_bat15;
reg [D*(LOC_BW-1)-1:0] loc_rdata_buff;
integer bi;
reg [4:0] loc_sram_buff_w0[0:255],loc_sram_buff_w1[0:255],loc_sram_buff_w2[0:255],loc_sram_buff_w3[0:255],loc_sram_buff_w4[0:255],loc_sram_buff_w5[0:255],loc_sram_buff_w6[0:255],loc_sram_buff_w7[0:255],loc_sram_buff_w8[0:255],loc_sram_buff_w9[0:255],loc_sram_buff_w10[0:255],loc_sram_buff_w11[0:255],loc_sram_buff_w12[0:255],loc_sram_buff_w13[0:255],loc_sram_buff_w14[0:255],loc_sram_buff_w15[0:255];
always @* begin 
	{loc_sram_buff_w0[0],loc_sram_buff_w0[1],loc_sram_buff_w0[2],loc_sram_buff_w0[3],loc_sram_buff_w0[4],loc_sram_buff_w0[5],loc_sram_buff_w0[6],loc_sram_buff_w0[7],loc_sram_buff_w0[8],loc_sram_buff_w0[9],loc_sram_buff_w0[10],loc_sram_buff_w0[11],loc_sram_buff_w0[12],loc_sram_buff_w0[13],loc_sram_buff_w0[14],loc_sram_buff_w0[15],loc_sram_buff_w0[16],loc_sram_buff_w0[17],loc_sram_buff_w0[18],loc_sram_buff_w0[19],loc_sram_buff_w0[20],loc_sram_buff_w0[21],loc_sram_buff_w0[22],loc_sram_buff_w0[23],loc_sram_buff_w0[24],loc_sram_buff_w0[25],loc_sram_buff_w0[26],loc_sram_buff_w0[27],loc_sram_buff_w0[28],loc_sram_buff_w0[29],loc_sram_buff_w0[30],loc_sram_buff_w0[31],loc_sram_buff_w0[32],loc_sram_buff_w0[33],loc_sram_buff_w0[34],loc_sram_buff_w0[35],loc_sram_buff_w0[36],loc_sram_buff_w0[37],loc_sram_buff_w0[38],loc_sram_buff_w0[39],loc_sram_buff_w0[40],loc_sram_buff_w0[41],loc_sram_buff_w0[42],loc_sram_buff_w0[43],loc_sram_buff_w0[44],loc_sram_buff_w0[45],loc_sram_buff_w0[46],loc_sram_buff_w0[47],loc_sram_buff_w0[48],loc_sram_buff_w0[49],loc_sram_buff_w0[50],loc_sram_buff_w0[51],loc_sram_buff_w0[52],loc_sram_buff_w0[53],loc_sram_buff_w0[54],loc_sram_buff_w0[55],loc_sram_buff_w0[56],loc_sram_buff_w0[57],loc_sram_buff_w0[58],loc_sram_buff_w0[59],loc_sram_buff_w0[60],loc_sram_buff_w0[61],loc_sram_buff_w0[62],loc_sram_buff_w0[63],loc_sram_buff_w0[64],loc_sram_buff_w0[65],loc_sram_buff_w0[66],loc_sram_buff_w0[67],loc_sram_buff_w0[68],loc_sram_buff_w0[69],loc_sram_buff_w0[70],loc_sram_buff_w0[71],loc_sram_buff_w0[72],loc_sram_buff_w0[73],loc_sram_buff_w0[74],loc_sram_buff_w0[75],loc_sram_buff_w0[76],loc_sram_buff_w0[77],loc_sram_buff_w0[78],loc_sram_buff_w0[79],loc_sram_buff_w0[80],loc_sram_buff_w0[81],loc_sram_buff_w0[82],loc_sram_buff_w0[83],loc_sram_buff_w0[84],loc_sram_buff_w0[85],loc_sram_buff_w0[86],loc_sram_buff_w0[87],loc_sram_buff_w0[88],loc_sram_buff_w0[89],loc_sram_buff_w0[90],loc_sram_buff_w0[91],loc_sram_buff_w0[92],loc_sram_buff_w0[93],loc_sram_buff_w0[94],loc_sram_buff_w0[95],loc_sram_buff_w0[96],loc_sram_buff_w0[97],loc_sram_buff_w0[98],loc_sram_buff_w0[99],loc_sram_buff_w0[100],loc_sram_buff_w0[101],loc_sram_buff_w0[102],loc_sram_buff_w0[103],loc_sram_buff_w0[104],loc_sram_buff_w0[105],loc_sram_buff_w0[106],loc_sram_buff_w0[107],loc_sram_buff_w0[108],loc_sram_buff_w0[109],loc_sram_buff_w0[110],loc_sram_buff_w0[111],loc_sram_buff_w0[112],loc_sram_buff_w0[113],loc_sram_buff_w0[114],loc_sram_buff_w0[115],loc_sram_buff_w0[116],loc_sram_buff_w0[117],loc_sram_buff_w0[118],loc_sram_buff_w0[119],loc_sram_buff_w0[120],loc_sram_buff_w0[121],loc_sram_buff_w0[122],loc_sram_buff_w0[123],loc_sram_buff_w0[124],loc_sram_buff_w0[125],loc_sram_buff_w0[126],loc_sram_buff_w0[127],loc_sram_buff_w0[128],loc_sram_buff_w0[129],loc_sram_buff_w0[130],loc_sram_buff_w0[131],loc_sram_buff_w0[132],loc_sram_buff_w0[133],loc_sram_buff_w0[134],loc_sram_buff_w0[135],loc_sram_buff_w0[136],loc_sram_buff_w0[137],loc_sram_buff_w0[138],loc_sram_buff_w0[139],loc_sram_buff_w0[140],loc_sram_buff_w0[141],loc_sram_buff_w0[142],loc_sram_buff_w0[143],loc_sram_buff_w0[144],loc_sram_buff_w0[145],loc_sram_buff_w0[146],loc_sram_buff_w0[147],loc_sram_buff_w0[148],loc_sram_buff_w0[149],loc_sram_buff_w0[150],loc_sram_buff_w0[151],loc_sram_buff_w0[152],loc_sram_buff_w0[153],loc_sram_buff_w0[154],loc_sram_buff_w0[155],loc_sram_buff_w0[156],loc_sram_buff_w0[157],loc_sram_buff_w0[158],loc_sram_buff_w0[159],loc_sram_buff_w0[160],loc_sram_buff_w0[161],loc_sram_buff_w0[162],loc_sram_buff_w0[163],loc_sram_buff_w0[164],loc_sram_buff_w0[165],loc_sram_buff_w0[166],loc_sram_buff_w0[167],loc_sram_buff_w0[168],loc_sram_buff_w0[169],loc_sram_buff_w0[170],loc_sram_buff_w0[171],loc_sram_buff_w0[172],loc_sram_buff_w0[173],loc_sram_buff_w0[174],loc_sram_buff_w0[175],loc_sram_buff_w0[176],loc_sram_buff_w0[177],loc_sram_buff_w0[178],loc_sram_buff_w0[179],loc_sram_buff_w0[180],loc_sram_buff_w0[181],loc_sram_buff_w0[182],loc_sram_buff_w0[183],loc_sram_buff_w0[184],loc_sram_buff_w0[185],loc_sram_buff_w0[186],loc_sram_buff_w0[187],loc_sram_buff_w0[188],loc_sram_buff_w0[189],loc_sram_buff_w0[190],loc_sram_buff_w0[191],loc_sram_buff_w0[192],loc_sram_buff_w0[193],loc_sram_buff_w0[194],loc_sram_buff_w0[195],loc_sram_buff_w0[196],loc_sram_buff_w0[197],loc_sram_buff_w0[198],loc_sram_buff_w0[199],loc_sram_buff_w0[200],loc_sram_buff_w0[201],loc_sram_buff_w0[202],loc_sram_buff_w0[203],loc_sram_buff_w0[204],loc_sram_buff_w0[205],loc_sram_buff_w0[206],loc_sram_buff_w0[207],loc_sram_buff_w0[208],loc_sram_buff_w0[209],loc_sram_buff_w0[210],loc_sram_buff_w0[211],loc_sram_buff_w0[212],loc_sram_buff_w0[213],loc_sram_buff_w0[214],loc_sram_buff_w0[215],loc_sram_buff_w0[216],loc_sram_buff_w0[217],loc_sram_buff_w0[218],loc_sram_buff_w0[219],loc_sram_buff_w0[220],loc_sram_buff_w0[221],loc_sram_buff_w0[222],loc_sram_buff_w0[223],loc_sram_buff_w0[224],loc_sram_buff_w0[225],loc_sram_buff_w0[226],loc_sram_buff_w0[227],loc_sram_buff_w0[228],loc_sram_buff_w0[229],loc_sram_buff_w0[230],loc_sram_buff_w0[231],loc_sram_buff_w0[232],loc_sram_buff_w0[233],loc_sram_buff_w0[234],loc_sram_buff_w0[235],loc_sram_buff_w0[236],loc_sram_buff_w0[237],loc_sram_buff_w0[238],loc_sram_buff_w0[239],loc_sram_buff_w0[240],loc_sram_buff_w0[241],loc_sram_buff_w0[242],loc_sram_buff_w0[243],loc_sram_buff_w0[244],loc_sram_buff_w0[245],loc_sram_buff_w0[246],loc_sram_buff_w0[247],loc_sram_buff_w0[248],loc_sram_buff_w0[249],loc_sram_buff_w0[250],loc_sram_buff_w0[251],loc_sram_buff_w0[252],loc_sram_buff_w0[253],loc_sram_buff_w0[254],loc_sram_buff_w0[255]} = loc_sram_rdata0;
	{loc_sram_buff_w1[0],loc_sram_buff_w1[1],loc_sram_buff_w1[2],loc_sram_buff_w1[3],loc_sram_buff_w1[4],loc_sram_buff_w1[5],loc_sram_buff_w1[6],loc_sram_buff_w1[7],loc_sram_buff_w1[8],loc_sram_buff_w1[9],loc_sram_buff_w1[10],loc_sram_buff_w1[11],loc_sram_buff_w1[12],loc_sram_buff_w1[13],loc_sram_buff_w1[14],loc_sram_buff_w1[15],loc_sram_buff_w1[16],loc_sram_buff_w1[17],loc_sram_buff_w1[18],loc_sram_buff_w1[19],loc_sram_buff_w1[20],loc_sram_buff_w1[21],loc_sram_buff_w1[22],loc_sram_buff_w1[23],loc_sram_buff_w1[24],loc_sram_buff_w1[25],loc_sram_buff_w1[26],loc_sram_buff_w1[27],loc_sram_buff_w1[28],loc_sram_buff_w1[29],loc_sram_buff_w1[30],loc_sram_buff_w1[31],loc_sram_buff_w1[32],loc_sram_buff_w1[33],loc_sram_buff_w1[34],loc_sram_buff_w1[35],loc_sram_buff_w1[36],loc_sram_buff_w1[37],loc_sram_buff_w1[38],loc_sram_buff_w1[39],loc_sram_buff_w1[40],loc_sram_buff_w1[41],loc_sram_buff_w1[42],loc_sram_buff_w1[43],loc_sram_buff_w1[44],loc_sram_buff_w1[45],loc_sram_buff_w1[46],loc_sram_buff_w1[47],loc_sram_buff_w1[48],loc_sram_buff_w1[49],loc_sram_buff_w1[50],loc_sram_buff_w1[51],loc_sram_buff_w1[52],loc_sram_buff_w1[53],loc_sram_buff_w1[54],loc_sram_buff_w1[55],loc_sram_buff_w1[56],loc_sram_buff_w1[57],loc_sram_buff_w1[58],loc_sram_buff_w1[59],loc_sram_buff_w1[60],loc_sram_buff_w1[61],loc_sram_buff_w1[62],loc_sram_buff_w1[63],loc_sram_buff_w1[64],loc_sram_buff_w1[65],loc_sram_buff_w1[66],loc_sram_buff_w1[67],loc_sram_buff_w1[68],loc_sram_buff_w1[69],loc_sram_buff_w1[70],loc_sram_buff_w1[71],loc_sram_buff_w1[72],loc_sram_buff_w1[73],loc_sram_buff_w1[74],loc_sram_buff_w1[75],loc_sram_buff_w1[76],loc_sram_buff_w1[77],loc_sram_buff_w1[78],loc_sram_buff_w1[79],loc_sram_buff_w1[80],loc_sram_buff_w1[81],loc_sram_buff_w1[82],loc_sram_buff_w1[83],loc_sram_buff_w1[84],loc_sram_buff_w1[85],loc_sram_buff_w1[86],loc_sram_buff_w1[87],loc_sram_buff_w1[88],loc_sram_buff_w1[89],loc_sram_buff_w1[90],loc_sram_buff_w1[91],loc_sram_buff_w1[92],loc_sram_buff_w1[93],loc_sram_buff_w1[94],loc_sram_buff_w1[95],loc_sram_buff_w1[96],loc_sram_buff_w1[97],loc_sram_buff_w1[98],loc_sram_buff_w1[99],loc_sram_buff_w1[100],loc_sram_buff_w1[101],loc_sram_buff_w1[102],loc_sram_buff_w1[103],loc_sram_buff_w1[104],loc_sram_buff_w1[105],loc_sram_buff_w1[106],loc_sram_buff_w1[107],loc_sram_buff_w1[108],loc_sram_buff_w1[109],loc_sram_buff_w1[110],loc_sram_buff_w1[111],loc_sram_buff_w1[112],loc_sram_buff_w1[113],loc_sram_buff_w1[114],loc_sram_buff_w1[115],loc_sram_buff_w1[116],loc_sram_buff_w1[117],loc_sram_buff_w1[118],loc_sram_buff_w1[119],loc_sram_buff_w1[120],loc_sram_buff_w1[121],loc_sram_buff_w1[122],loc_sram_buff_w1[123],loc_sram_buff_w1[124],loc_sram_buff_w1[125],loc_sram_buff_w1[126],loc_sram_buff_w1[127],loc_sram_buff_w1[128],loc_sram_buff_w1[129],loc_sram_buff_w1[130],loc_sram_buff_w1[131],loc_sram_buff_w1[132],loc_sram_buff_w1[133],loc_sram_buff_w1[134],loc_sram_buff_w1[135],loc_sram_buff_w1[136],loc_sram_buff_w1[137],loc_sram_buff_w1[138],loc_sram_buff_w1[139],loc_sram_buff_w1[140],loc_sram_buff_w1[141],loc_sram_buff_w1[142],loc_sram_buff_w1[143],loc_sram_buff_w1[144],loc_sram_buff_w1[145],loc_sram_buff_w1[146],loc_sram_buff_w1[147],loc_sram_buff_w1[148],loc_sram_buff_w1[149],loc_sram_buff_w1[150],loc_sram_buff_w1[151],loc_sram_buff_w1[152],loc_sram_buff_w1[153],loc_sram_buff_w1[154],loc_sram_buff_w1[155],loc_sram_buff_w1[156],loc_sram_buff_w1[157],loc_sram_buff_w1[158],loc_sram_buff_w1[159],loc_sram_buff_w1[160],loc_sram_buff_w1[161],loc_sram_buff_w1[162],loc_sram_buff_w1[163],loc_sram_buff_w1[164],loc_sram_buff_w1[165],loc_sram_buff_w1[166],loc_sram_buff_w1[167],loc_sram_buff_w1[168],loc_sram_buff_w1[169],loc_sram_buff_w1[170],loc_sram_buff_w1[171],loc_sram_buff_w1[172],loc_sram_buff_w1[173],loc_sram_buff_w1[174],loc_sram_buff_w1[175],loc_sram_buff_w1[176],loc_sram_buff_w1[177],loc_sram_buff_w1[178],loc_sram_buff_w1[179],loc_sram_buff_w1[180],loc_sram_buff_w1[181],loc_sram_buff_w1[182],loc_sram_buff_w1[183],loc_sram_buff_w1[184],loc_sram_buff_w1[185],loc_sram_buff_w1[186],loc_sram_buff_w1[187],loc_sram_buff_w1[188],loc_sram_buff_w1[189],loc_sram_buff_w1[190],loc_sram_buff_w1[191],loc_sram_buff_w1[192],loc_sram_buff_w1[193],loc_sram_buff_w1[194],loc_sram_buff_w1[195],loc_sram_buff_w1[196],loc_sram_buff_w1[197],loc_sram_buff_w1[198],loc_sram_buff_w1[199],loc_sram_buff_w1[200],loc_sram_buff_w1[201],loc_sram_buff_w1[202],loc_sram_buff_w1[203],loc_sram_buff_w1[204],loc_sram_buff_w1[205],loc_sram_buff_w1[206],loc_sram_buff_w1[207],loc_sram_buff_w1[208],loc_sram_buff_w1[209],loc_sram_buff_w1[210],loc_sram_buff_w1[211],loc_sram_buff_w1[212],loc_sram_buff_w1[213],loc_sram_buff_w1[214],loc_sram_buff_w1[215],loc_sram_buff_w1[216],loc_sram_buff_w1[217],loc_sram_buff_w1[218],loc_sram_buff_w1[219],loc_sram_buff_w1[220],loc_sram_buff_w1[221],loc_sram_buff_w1[222],loc_sram_buff_w1[223],loc_sram_buff_w1[224],loc_sram_buff_w1[225],loc_sram_buff_w1[226],loc_sram_buff_w1[227],loc_sram_buff_w1[228],loc_sram_buff_w1[229],loc_sram_buff_w1[230],loc_sram_buff_w1[231],loc_sram_buff_w1[232],loc_sram_buff_w1[233],loc_sram_buff_w1[234],loc_sram_buff_w1[235],loc_sram_buff_w1[236],loc_sram_buff_w1[237],loc_sram_buff_w1[238],loc_sram_buff_w1[239],loc_sram_buff_w1[240],loc_sram_buff_w1[241],loc_sram_buff_w1[242],loc_sram_buff_w1[243],loc_sram_buff_w1[244],loc_sram_buff_w1[245],loc_sram_buff_w1[246],loc_sram_buff_w1[247],loc_sram_buff_w1[248],loc_sram_buff_w1[249],loc_sram_buff_w1[250],loc_sram_buff_w1[251],loc_sram_buff_w1[252],loc_sram_buff_w1[253],loc_sram_buff_w1[254],loc_sram_buff_w1[255]} = loc_sram_rdata1;
	{loc_sram_buff_w2[0],loc_sram_buff_w2[1],loc_sram_buff_w2[2],loc_sram_buff_w2[3],loc_sram_buff_w2[4],loc_sram_buff_w2[5],loc_sram_buff_w2[6],loc_sram_buff_w2[7],loc_sram_buff_w2[8],loc_sram_buff_w2[9],loc_sram_buff_w2[10],loc_sram_buff_w2[11],loc_sram_buff_w2[12],loc_sram_buff_w2[13],loc_sram_buff_w2[14],loc_sram_buff_w2[15],loc_sram_buff_w2[16],loc_sram_buff_w2[17],loc_sram_buff_w2[18],loc_sram_buff_w2[19],loc_sram_buff_w2[20],loc_sram_buff_w2[21],loc_sram_buff_w2[22],loc_sram_buff_w2[23],loc_sram_buff_w2[24],loc_sram_buff_w2[25],loc_sram_buff_w2[26],loc_sram_buff_w2[27],loc_sram_buff_w2[28],loc_sram_buff_w2[29],loc_sram_buff_w2[30],loc_sram_buff_w2[31],loc_sram_buff_w2[32],loc_sram_buff_w2[33],loc_sram_buff_w2[34],loc_sram_buff_w2[35],loc_sram_buff_w2[36],loc_sram_buff_w2[37],loc_sram_buff_w2[38],loc_sram_buff_w2[39],loc_sram_buff_w2[40],loc_sram_buff_w2[41],loc_sram_buff_w2[42],loc_sram_buff_w2[43],loc_sram_buff_w2[44],loc_sram_buff_w2[45],loc_sram_buff_w2[46],loc_sram_buff_w2[47],loc_sram_buff_w2[48],loc_sram_buff_w2[49],loc_sram_buff_w2[50],loc_sram_buff_w2[51],loc_sram_buff_w2[52],loc_sram_buff_w2[53],loc_sram_buff_w2[54],loc_sram_buff_w2[55],loc_sram_buff_w2[56],loc_sram_buff_w2[57],loc_sram_buff_w2[58],loc_sram_buff_w2[59],loc_sram_buff_w2[60],loc_sram_buff_w2[61],loc_sram_buff_w2[62],loc_sram_buff_w2[63],loc_sram_buff_w2[64],loc_sram_buff_w2[65],loc_sram_buff_w2[66],loc_sram_buff_w2[67],loc_sram_buff_w2[68],loc_sram_buff_w2[69],loc_sram_buff_w2[70],loc_sram_buff_w2[71],loc_sram_buff_w2[72],loc_sram_buff_w2[73],loc_sram_buff_w2[74],loc_sram_buff_w2[75],loc_sram_buff_w2[76],loc_sram_buff_w2[77],loc_sram_buff_w2[78],loc_sram_buff_w2[79],loc_sram_buff_w2[80],loc_sram_buff_w2[81],loc_sram_buff_w2[82],loc_sram_buff_w2[83],loc_sram_buff_w2[84],loc_sram_buff_w2[85],loc_sram_buff_w2[86],loc_sram_buff_w2[87],loc_sram_buff_w2[88],loc_sram_buff_w2[89],loc_sram_buff_w2[90],loc_sram_buff_w2[91],loc_sram_buff_w2[92],loc_sram_buff_w2[93],loc_sram_buff_w2[94],loc_sram_buff_w2[95],loc_sram_buff_w2[96],loc_sram_buff_w2[97],loc_sram_buff_w2[98],loc_sram_buff_w2[99],loc_sram_buff_w2[100],loc_sram_buff_w2[101],loc_sram_buff_w2[102],loc_sram_buff_w2[103],loc_sram_buff_w2[104],loc_sram_buff_w2[105],loc_sram_buff_w2[106],loc_sram_buff_w2[107],loc_sram_buff_w2[108],loc_sram_buff_w2[109],loc_sram_buff_w2[110],loc_sram_buff_w2[111],loc_sram_buff_w2[112],loc_sram_buff_w2[113],loc_sram_buff_w2[114],loc_sram_buff_w2[115],loc_sram_buff_w2[116],loc_sram_buff_w2[117],loc_sram_buff_w2[118],loc_sram_buff_w2[119],loc_sram_buff_w2[120],loc_sram_buff_w2[121],loc_sram_buff_w2[122],loc_sram_buff_w2[123],loc_sram_buff_w2[124],loc_sram_buff_w2[125],loc_sram_buff_w2[126],loc_sram_buff_w2[127],loc_sram_buff_w2[128],loc_sram_buff_w2[129],loc_sram_buff_w2[130],loc_sram_buff_w2[131],loc_sram_buff_w2[132],loc_sram_buff_w2[133],loc_sram_buff_w2[134],loc_sram_buff_w2[135],loc_sram_buff_w2[136],loc_sram_buff_w2[137],loc_sram_buff_w2[138],loc_sram_buff_w2[139],loc_sram_buff_w2[140],loc_sram_buff_w2[141],loc_sram_buff_w2[142],loc_sram_buff_w2[143],loc_sram_buff_w2[144],loc_sram_buff_w2[145],loc_sram_buff_w2[146],loc_sram_buff_w2[147],loc_sram_buff_w2[148],loc_sram_buff_w2[149],loc_sram_buff_w2[150],loc_sram_buff_w2[151],loc_sram_buff_w2[152],loc_sram_buff_w2[153],loc_sram_buff_w2[154],loc_sram_buff_w2[155],loc_sram_buff_w2[156],loc_sram_buff_w2[157],loc_sram_buff_w2[158],loc_sram_buff_w2[159],loc_sram_buff_w2[160],loc_sram_buff_w2[161],loc_sram_buff_w2[162],loc_sram_buff_w2[163],loc_sram_buff_w2[164],loc_sram_buff_w2[165],loc_sram_buff_w2[166],loc_sram_buff_w2[167],loc_sram_buff_w2[168],loc_sram_buff_w2[169],loc_sram_buff_w2[170],loc_sram_buff_w2[171],loc_sram_buff_w2[172],loc_sram_buff_w2[173],loc_sram_buff_w2[174],loc_sram_buff_w2[175],loc_sram_buff_w2[176],loc_sram_buff_w2[177],loc_sram_buff_w2[178],loc_sram_buff_w2[179],loc_sram_buff_w2[180],loc_sram_buff_w2[181],loc_sram_buff_w2[182],loc_sram_buff_w2[183],loc_sram_buff_w2[184],loc_sram_buff_w2[185],loc_sram_buff_w2[186],loc_sram_buff_w2[187],loc_sram_buff_w2[188],loc_sram_buff_w2[189],loc_sram_buff_w2[190],loc_sram_buff_w2[191],loc_sram_buff_w2[192],loc_sram_buff_w2[193],loc_sram_buff_w2[194],loc_sram_buff_w2[195],loc_sram_buff_w2[196],loc_sram_buff_w2[197],loc_sram_buff_w2[198],loc_sram_buff_w2[199],loc_sram_buff_w2[200],loc_sram_buff_w2[201],loc_sram_buff_w2[202],loc_sram_buff_w2[203],loc_sram_buff_w2[204],loc_sram_buff_w2[205],loc_sram_buff_w2[206],loc_sram_buff_w2[207],loc_sram_buff_w2[208],loc_sram_buff_w2[209],loc_sram_buff_w2[210],loc_sram_buff_w2[211],loc_sram_buff_w2[212],loc_sram_buff_w2[213],loc_sram_buff_w2[214],loc_sram_buff_w2[215],loc_sram_buff_w2[216],loc_sram_buff_w2[217],loc_sram_buff_w2[218],loc_sram_buff_w2[219],loc_sram_buff_w2[220],loc_sram_buff_w2[221],loc_sram_buff_w2[222],loc_sram_buff_w2[223],loc_sram_buff_w2[224],loc_sram_buff_w2[225],loc_sram_buff_w2[226],loc_sram_buff_w2[227],loc_sram_buff_w2[228],loc_sram_buff_w2[229],loc_sram_buff_w2[230],loc_sram_buff_w2[231],loc_sram_buff_w2[232],loc_sram_buff_w2[233],loc_sram_buff_w2[234],loc_sram_buff_w2[235],loc_sram_buff_w2[236],loc_sram_buff_w2[237],loc_sram_buff_w2[238],loc_sram_buff_w2[239],loc_sram_buff_w2[240],loc_sram_buff_w2[241],loc_sram_buff_w2[242],loc_sram_buff_w2[243],loc_sram_buff_w2[244],loc_sram_buff_w2[245],loc_sram_buff_w2[246],loc_sram_buff_w2[247],loc_sram_buff_w2[248],loc_sram_buff_w2[249],loc_sram_buff_w2[250],loc_sram_buff_w2[251],loc_sram_buff_w2[252],loc_sram_buff_w2[253],loc_sram_buff_w2[254],loc_sram_buff_w2[255]} = loc_sram_rdata2;
	{loc_sram_buff_w3[0],loc_sram_buff_w3[1],loc_sram_buff_w3[2],loc_sram_buff_w3[3],loc_sram_buff_w3[4],loc_sram_buff_w3[5],loc_sram_buff_w3[6],loc_sram_buff_w3[7],loc_sram_buff_w3[8],loc_sram_buff_w3[9],loc_sram_buff_w3[10],loc_sram_buff_w3[11],loc_sram_buff_w3[12],loc_sram_buff_w3[13],loc_sram_buff_w3[14],loc_sram_buff_w3[15],loc_sram_buff_w3[16],loc_sram_buff_w3[17],loc_sram_buff_w3[18],loc_sram_buff_w3[19],loc_sram_buff_w3[20],loc_sram_buff_w3[21],loc_sram_buff_w3[22],loc_sram_buff_w3[23],loc_sram_buff_w3[24],loc_sram_buff_w3[25],loc_sram_buff_w3[26],loc_sram_buff_w3[27],loc_sram_buff_w3[28],loc_sram_buff_w3[29],loc_sram_buff_w3[30],loc_sram_buff_w3[31],loc_sram_buff_w3[32],loc_sram_buff_w3[33],loc_sram_buff_w3[34],loc_sram_buff_w3[35],loc_sram_buff_w3[36],loc_sram_buff_w3[37],loc_sram_buff_w3[38],loc_sram_buff_w3[39],loc_sram_buff_w3[40],loc_sram_buff_w3[41],loc_sram_buff_w3[42],loc_sram_buff_w3[43],loc_sram_buff_w3[44],loc_sram_buff_w3[45],loc_sram_buff_w3[46],loc_sram_buff_w3[47],loc_sram_buff_w3[48],loc_sram_buff_w3[49],loc_sram_buff_w3[50],loc_sram_buff_w3[51],loc_sram_buff_w3[52],loc_sram_buff_w3[53],loc_sram_buff_w3[54],loc_sram_buff_w3[55],loc_sram_buff_w3[56],loc_sram_buff_w3[57],loc_sram_buff_w3[58],loc_sram_buff_w3[59],loc_sram_buff_w3[60],loc_sram_buff_w3[61],loc_sram_buff_w3[62],loc_sram_buff_w3[63],loc_sram_buff_w3[64],loc_sram_buff_w3[65],loc_sram_buff_w3[66],loc_sram_buff_w3[67],loc_sram_buff_w3[68],loc_sram_buff_w3[69],loc_sram_buff_w3[70],loc_sram_buff_w3[71],loc_sram_buff_w3[72],loc_sram_buff_w3[73],loc_sram_buff_w3[74],loc_sram_buff_w3[75],loc_sram_buff_w3[76],loc_sram_buff_w3[77],loc_sram_buff_w3[78],loc_sram_buff_w3[79],loc_sram_buff_w3[80],loc_sram_buff_w3[81],loc_sram_buff_w3[82],loc_sram_buff_w3[83],loc_sram_buff_w3[84],loc_sram_buff_w3[85],loc_sram_buff_w3[86],loc_sram_buff_w3[87],loc_sram_buff_w3[88],loc_sram_buff_w3[89],loc_sram_buff_w3[90],loc_sram_buff_w3[91],loc_sram_buff_w3[92],loc_sram_buff_w3[93],loc_sram_buff_w3[94],loc_sram_buff_w3[95],loc_sram_buff_w3[96],loc_sram_buff_w3[97],loc_sram_buff_w3[98],loc_sram_buff_w3[99],loc_sram_buff_w3[100],loc_sram_buff_w3[101],loc_sram_buff_w3[102],loc_sram_buff_w3[103],loc_sram_buff_w3[104],loc_sram_buff_w3[105],loc_sram_buff_w3[106],loc_sram_buff_w3[107],loc_sram_buff_w3[108],loc_sram_buff_w3[109],loc_sram_buff_w3[110],loc_sram_buff_w3[111],loc_sram_buff_w3[112],loc_sram_buff_w3[113],loc_sram_buff_w3[114],loc_sram_buff_w3[115],loc_sram_buff_w3[116],loc_sram_buff_w3[117],loc_sram_buff_w3[118],loc_sram_buff_w3[119],loc_sram_buff_w3[120],loc_sram_buff_w3[121],loc_sram_buff_w3[122],loc_sram_buff_w3[123],loc_sram_buff_w3[124],loc_sram_buff_w3[125],loc_sram_buff_w3[126],loc_sram_buff_w3[127],loc_sram_buff_w3[128],loc_sram_buff_w3[129],loc_sram_buff_w3[130],loc_sram_buff_w3[131],loc_sram_buff_w3[132],loc_sram_buff_w3[133],loc_sram_buff_w3[134],loc_sram_buff_w3[135],loc_sram_buff_w3[136],loc_sram_buff_w3[137],loc_sram_buff_w3[138],loc_sram_buff_w3[139],loc_sram_buff_w3[140],loc_sram_buff_w3[141],loc_sram_buff_w3[142],loc_sram_buff_w3[143],loc_sram_buff_w3[144],loc_sram_buff_w3[145],loc_sram_buff_w3[146],loc_sram_buff_w3[147],loc_sram_buff_w3[148],loc_sram_buff_w3[149],loc_sram_buff_w3[150],loc_sram_buff_w3[151],loc_sram_buff_w3[152],loc_sram_buff_w3[153],loc_sram_buff_w3[154],loc_sram_buff_w3[155],loc_sram_buff_w3[156],loc_sram_buff_w3[157],loc_sram_buff_w3[158],loc_sram_buff_w3[159],loc_sram_buff_w3[160],loc_sram_buff_w3[161],loc_sram_buff_w3[162],loc_sram_buff_w3[163],loc_sram_buff_w3[164],loc_sram_buff_w3[165],loc_sram_buff_w3[166],loc_sram_buff_w3[167],loc_sram_buff_w3[168],loc_sram_buff_w3[169],loc_sram_buff_w3[170],loc_sram_buff_w3[171],loc_sram_buff_w3[172],loc_sram_buff_w3[173],loc_sram_buff_w3[174],loc_sram_buff_w3[175],loc_sram_buff_w3[176],loc_sram_buff_w3[177],loc_sram_buff_w3[178],loc_sram_buff_w3[179],loc_sram_buff_w3[180],loc_sram_buff_w3[181],loc_sram_buff_w3[182],loc_sram_buff_w3[183],loc_sram_buff_w3[184],loc_sram_buff_w3[185],loc_sram_buff_w3[186],loc_sram_buff_w3[187],loc_sram_buff_w3[188],loc_sram_buff_w3[189],loc_sram_buff_w3[190],loc_sram_buff_w3[191],loc_sram_buff_w3[192],loc_sram_buff_w3[193],loc_sram_buff_w3[194],loc_sram_buff_w3[195],loc_sram_buff_w3[196],loc_sram_buff_w3[197],loc_sram_buff_w3[198],loc_sram_buff_w3[199],loc_sram_buff_w3[200],loc_sram_buff_w3[201],loc_sram_buff_w3[202],loc_sram_buff_w3[203],loc_sram_buff_w3[204],loc_sram_buff_w3[205],loc_sram_buff_w3[206],loc_sram_buff_w3[207],loc_sram_buff_w3[208],loc_sram_buff_w3[209],loc_sram_buff_w3[210],loc_sram_buff_w3[211],loc_sram_buff_w3[212],loc_sram_buff_w3[213],loc_sram_buff_w3[214],loc_sram_buff_w3[215],loc_sram_buff_w3[216],loc_sram_buff_w3[217],loc_sram_buff_w3[218],loc_sram_buff_w3[219],loc_sram_buff_w3[220],loc_sram_buff_w3[221],loc_sram_buff_w3[222],loc_sram_buff_w3[223],loc_sram_buff_w3[224],loc_sram_buff_w3[225],loc_sram_buff_w3[226],loc_sram_buff_w3[227],loc_sram_buff_w3[228],loc_sram_buff_w3[229],loc_sram_buff_w3[230],loc_sram_buff_w3[231],loc_sram_buff_w3[232],loc_sram_buff_w3[233],loc_sram_buff_w3[234],loc_sram_buff_w3[235],loc_sram_buff_w3[236],loc_sram_buff_w3[237],loc_sram_buff_w3[238],loc_sram_buff_w3[239],loc_sram_buff_w3[240],loc_sram_buff_w3[241],loc_sram_buff_w3[242],loc_sram_buff_w3[243],loc_sram_buff_w3[244],loc_sram_buff_w3[245],loc_sram_buff_w3[246],loc_sram_buff_w3[247],loc_sram_buff_w3[248],loc_sram_buff_w3[249],loc_sram_buff_w3[250],loc_sram_buff_w3[251],loc_sram_buff_w3[252],loc_sram_buff_w3[253],loc_sram_buff_w3[254],loc_sram_buff_w3[255]} = loc_sram_rdata3;
	{loc_sram_buff_w4[0],loc_sram_buff_w4[1],loc_sram_buff_w4[2],loc_sram_buff_w4[3],loc_sram_buff_w4[4],loc_sram_buff_w4[5],loc_sram_buff_w4[6],loc_sram_buff_w4[7],loc_sram_buff_w4[8],loc_sram_buff_w4[9],loc_sram_buff_w4[10],loc_sram_buff_w4[11],loc_sram_buff_w4[12],loc_sram_buff_w4[13],loc_sram_buff_w4[14],loc_sram_buff_w4[15],loc_sram_buff_w4[16],loc_sram_buff_w4[17],loc_sram_buff_w4[18],loc_sram_buff_w4[19],loc_sram_buff_w4[20],loc_sram_buff_w4[21],loc_sram_buff_w4[22],loc_sram_buff_w4[23],loc_sram_buff_w4[24],loc_sram_buff_w4[25],loc_sram_buff_w4[26],loc_sram_buff_w4[27],loc_sram_buff_w4[28],loc_sram_buff_w4[29],loc_sram_buff_w4[30],loc_sram_buff_w4[31],loc_sram_buff_w4[32],loc_sram_buff_w4[33],loc_sram_buff_w4[34],loc_sram_buff_w4[35],loc_sram_buff_w4[36],loc_sram_buff_w4[37],loc_sram_buff_w4[38],loc_sram_buff_w4[39],loc_sram_buff_w4[40],loc_sram_buff_w4[41],loc_sram_buff_w4[42],loc_sram_buff_w4[43],loc_sram_buff_w4[44],loc_sram_buff_w4[45],loc_sram_buff_w4[46],loc_sram_buff_w4[47],loc_sram_buff_w4[48],loc_sram_buff_w4[49],loc_sram_buff_w4[50],loc_sram_buff_w4[51],loc_sram_buff_w4[52],loc_sram_buff_w4[53],loc_sram_buff_w4[54],loc_sram_buff_w4[55],loc_sram_buff_w4[56],loc_sram_buff_w4[57],loc_sram_buff_w4[58],loc_sram_buff_w4[59],loc_sram_buff_w4[60],loc_sram_buff_w4[61],loc_sram_buff_w4[62],loc_sram_buff_w4[63],loc_sram_buff_w4[64],loc_sram_buff_w4[65],loc_sram_buff_w4[66],loc_sram_buff_w4[67],loc_sram_buff_w4[68],loc_sram_buff_w4[69],loc_sram_buff_w4[70],loc_sram_buff_w4[71],loc_sram_buff_w4[72],loc_sram_buff_w4[73],loc_sram_buff_w4[74],loc_sram_buff_w4[75],loc_sram_buff_w4[76],loc_sram_buff_w4[77],loc_sram_buff_w4[78],loc_sram_buff_w4[79],loc_sram_buff_w4[80],loc_sram_buff_w4[81],loc_sram_buff_w4[82],loc_sram_buff_w4[83],loc_sram_buff_w4[84],loc_sram_buff_w4[85],loc_sram_buff_w4[86],loc_sram_buff_w4[87],loc_sram_buff_w4[88],loc_sram_buff_w4[89],loc_sram_buff_w4[90],loc_sram_buff_w4[91],loc_sram_buff_w4[92],loc_sram_buff_w4[93],loc_sram_buff_w4[94],loc_sram_buff_w4[95],loc_sram_buff_w4[96],loc_sram_buff_w4[97],loc_sram_buff_w4[98],loc_sram_buff_w4[99],loc_sram_buff_w4[100],loc_sram_buff_w4[101],loc_sram_buff_w4[102],loc_sram_buff_w4[103],loc_sram_buff_w4[104],loc_sram_buff_w4[105],loc_sram_buff_w4[106],loc_sram_buff_w4[107],loc_sram_buff_w4[108],loc_sram_buff_w4[109],loc_sram_buff_w4[110],loc_sram_buff_w4[111],loc_sram_buff_w4[112],loc_sram_buff_w4[113],loc_sram_buff_w4[114],loc_sram_buff_w4[115],loc_sram_buff_w4[116],loc_sram_buff_w4[117],loc_sram_buff_w4[118],loc_sram_buff_w4[119],loc_sram_buff_w4[120],loc_sram_buff_w4[121],loc_sram_buff_w4[122],loc_sram_buff_w4[123],loc_sram_buff_w4[124],loc_sram_buff_w4[125],loc_sram_buff_w4[126],loc_sram_buff_w4[127],loc_sram_buff_w4[128],loc_sram_buff_w4[129],loc_sram_buff_w4[130],loc_sram_buff_w4[131],loc_sram_buff_w4[132],loc_sram_buff_w4[133],loc_sram_buff_w4[134],loc_sram_buff_w4[135],loc_sram_buff_w4[136],loc_sram_buff_w4[137],loc_sram_buff_w4[138],loc_sram_buff_w4[139],loc_sram_buff_w4[140],loc_sram_buff_w4[141],loc_sram_buff_w4[142],loc_sram_buff_w4[143],loc_sram_buff_w4[144],loc_sram_buff_w4[145],loc_sram_buff_w4[146],loc_sram_buff_w4[147],loc_sram_buff_w4[148],loc_sram_buff_w4[149],loc_sram_buff_w4[150],loc_sram_buff_w4[151],loc_sram_buff_w4[152],loc_sram_buff_w4[153],loc_sram_buff_w4[154],loc_sram_buff_w4[155],loc_sram_buff_w4[156],loc_sram_buff_w4[157],loc_sram_buff_w4[158],loc_sram_buff_w4[159],loc_sram_buff_w4[160],loc_sram_buff_w4[161],loc_sram_buff_w4[162],loc_sram_buff_w4[163],loc_sram_buff_w4[164],loc_sram_buff_w4[165],loc_sram_buff_w4[166],loc_sram_buff_w4[167],loc_sram_buff_w4[168],loc_sram_buff_w4[169],loc_sram_buff_w4[170],loc_sram_buff_w4[171],loc_sram_buff_w4[172],loc_sram_buff_w4[173],loc_sram_buff_w4[174],loc_sram_buff_w4[175],loc_sram_buff_w4[176],loc_sram_buff_w4[177],loc_sram_buff_w4[178],loc_sram_buff_w4[179],loc_sram_buff_w4[180],loc_sram_buff_w4[181],loc_sram_buff_w4[182],loc_sram_buff_w4[183],loc_sram_buff_w4[184],loc_sram_buff_w4[185],loc_sram_buff_w4[186],loc_sram_buff_w4[187],loc_sram_buff_w4[188],loc_sram_buff_w4[189],loc_sram_buff_w4[190],loc_sram_buff_w4[191],loc_sram_buff_w4[192],loc_sram_buff_w4[193],loc_sram_buff_w4[194],loc_sram_buff_w4[195],loc_sram_buff_w4[196],loc_sram_buff_w4[197],loc_sram_buff_w4[198],loc_sram_buff_w4[199],loc_sram_buff_w4[200],loc_sram_buff_w4[201],loc_sram_buff_w4[202],loc_sram_buff_w4[203],loc_sram_buff_w4[204],loc_sram_buff_w4[205],loc_sram_buff_w4[206],loc_sram_buff_w4[207],loc_sram_buff_w4[208],loc_sram_buff_w4[209],loc_sram_buff_w4[210],loc_sram_buff_w4[211],loc_sram_buff_w4[212],loc_sram_buff_w4[213],loc_sram_buff_w4[214],loc_sram_buff_w4[215],loc_sram_buff_w4[216],loc_sram_buff_w4[217],loc_sram_buff_w4[218],loc_sram_buff_w4[219],loc_sram_buff_w4[220],loc_sram_buff_w4[221],loc_sram_buff_w4[222],loc_sram_buff_w4[223],loc_sram_buff_w4[224],loc_sram_buff_w4[225],loc_sram_buff_w4[226],loc_sram_buff_w4[227],loc_sram_buff_w4[228],loc_sram_buff_w4[229],loc_sram_buff_w4[230],loc_sram_buff_w4[231],loc_sram_buff_w4[232],loc_sram_buff_w4[233],loc_sram_buff_w4[234],loc_sram_buff_w4[235],loc_sram_buff_w4[236],loc_sram_buff_w4[237],loc_sram_buff_w4[238],loc_sram_buff_w4[239],loc_sram_buff_w4[240],loc_sram_buff_w4[241],loc_sram_buff_w4[242],loc_sram_buff_w4[243],loc_sram_buff_w4[244],loc_sram_buff_w4[245],loc_sram_buff_w4[246],loc_sram_buff_w4[247],loc_sram_buff_w4[248],loc_sram_buff_w4[249],loc_sram_buff_w4[250],loc_sram_buff_w4[251],loc_sram_buff_w4[252],loc_sram_buff_w4[253],loc_sram_buff_w4[254],loc_sram_buff_w4[255]} = loc_sram_rdata4;
	{loc_sram_buff_w5[0],loc_sram_buff_w5[1],loc_sram_buff_w5[2],loc_sram_buff_w5[3],loc_sram_buff_w5[4],loc_sram_buff_w5[5],loc_sram_buff_w5[6],loc_sram_buff_w5[7],loc_sram_buff_w5[8],loc_sram_buff_w5[9],loc_sram_buff_w5[10],loc_sram_buff_w5[11],loc_sram_buff_w5[12],loc_sram_buff_w5[13],loc_sram_buff_w5[14],loc_sram_buff_w5[15],loc_sram_buff_w5[16],loc_sram_buff_w5[17],loc_sram_buff_w5[18],loc_sram_buff_w5[19],loc_sram_buff_w5[20],loc_sram_buff_w5[21],loc_sram_buff_w5[22],loc_sram_buff_w5[23],loc_sram_buff_w5[24],loc_sram_buff_w5[25],loc_sram_buff_w5[26],loc_sram_buff_w5[27],loc_sram_buff_w5[28],loc_sram_buff_w5[29],loc_sram_buff_w5[30],loc_sram_buff_w5[31],loc_sram_buff_w5[32],loc_sram_buff_w5[33],loc_sram_buff_w5[34],loc_sram_buff_w5[35],loc_sram_buff_w5[36],loc_sram_buff_w5[37],loc_sram_buff_w5[38],loc_sram_buff_w5[39],loc_sram_buff_w5[40],loc_sram_buff_w5[41],loc_sram_buff_w5[42],loc_sram_buff_w5[43],loc_sram_buff_w5[44],loc_sram_buff_w5[45],loc_sram_buff_w5[46],loc_sram_buff_w5[47],loc_sram_buff_w5[48],loc_sram_buff_w5[49],loc_sram_buff_w5[50],loc_sram_buff_w5[51],loc_sram_buff_w5[52],loc_sram_buff_w5[53],loc_sram_buff_w5[54],loc_sram_buff_w5[55],loc_sram_buff_w5[56],loc_sram_buff_w5[57],loc_sram_buff_w5[58],loc_sram_buff_w5[59],loc_sram_buff_w5[60],loc_sram_buff_w5[61],loc_sram_buff_w5[62],loc_sram_buff_w5[63],loc_sram_buff_w5[64],loc_sram_buff_w5[65],loc_sram_buff_w5[66],loc_sram_buff_w5[67],loc_sram_buff_w5[68],loc_sram_buff_w5[69],loc_sram_buff_w5[70],loc_sram_buff_w5[71],loc_sram_buff_w5[72],loc_sram_buff_w5[73],loc_sram_buff_w5[74],loc_sram_buff_w5[75],loc_sram_buff_w5[76],loc_sram_buff_w5[77],loc_sram_buff_w5[78],loc_sram_buff_w5[79],loc_sram_buff_w5[80],loc_sram_buff_w5[81],loc_sram_buff_w5[82],loc_sram_buff_w5[83],loc_sram_buff_w5[84],loc_sram_buff_w5[85],loc_sram_buff_w5[86],loc_sram_buff_w5[87],loc_sram_buff_w5[88],loc_sram_buff_w5[89],loc_sram_buff_w5[90],loc_sram_buff_w5[91],loc_sram_buff_w5[92],loc_sram_buff_w5[93],loc_sram_buff_w5[94],loc_sram_buff_w5[95],loc_sram_buff_w5[96],loc_sram_buff_w5[97],loc_sram_buff_w5[98],loc_sram_buff_w5[99],loc_sram_buff_w5[100],loc_sram_buff_w5[101],loc_sram_buff_w5[102],loc_sram_buff_w5[103],loc_sram_buff_w5[104],loc_sram_buff_w5[105],loc_sram_buff_w5[106],loc_sram_buff_w5[107],loc_sram_buff_w5[108],loc_sram_buff_w5[109],loc_sram_buff_w5[110],loc_sram_buff_w5[111],loc_sram_buff_w5[112],loc_sram_buff_w5[113],loc_sram_buff_w5[114],loc_sram_buff_w5[115],loc_sram_buff_w5[116],loc_sram_buff_w5[117],loc_sram_buff_w5[118],loc_sram_buff_w5[119],loc_sram_buff_w5[120],loc_sram_buff_w5[121],loc_sram_buff_w5[122],loc_sram_buff_w5[123],loc_sram_buff_w5[124],loc_sram_buff_w5[125],loc_sram_buff_w5[126],loc_sram_buff_w5[127],loc_sram_buff_w5[128],loc_sram_buff_w5[129],loc_sram_buff_w5[130],loc_sram_buff_w5[131],loc_sram_buff_w5[132],loc_sram_buff_w5[133],loc_sram_buff_w5[134],loc_sram_buff_w5[135],loc_sram_buff_w5[136],loc_sram_buff_w5[137],loc_sram_buff_w5[138],loc_sram_buff_w5[139],loc_sram_buff_w5[140],loc_sram_buff_w5[141],loc_sram_buff_w5[142],loc_sram_buff_w5[143],loc_sram_buff_w5[144],loc_sram_buff_w5[145],loc_sram_buff_w5[146],loc_sram_buff_w5[147],loc_sram_buff_w5[148],loc_sram_buff_w5[149],loc_sram_buff_w5[150],loc_sram_buff_w5[151],loc_sram_buff_w5[152],loc_sram_buff_w5[153],loc_sram_buff_w5[154],loc_sram_buff_w5[155],loc_sram_buff_w5[156],loc_sram_buff_w5[157],loc_sram_buff_w5[158],loc_sram_buff_w5[159],loc_sram_buff_w5[160],loc_sram_buff_w5[161],loc_sram_buff_w5[162],loc_sram_buff_w5[163],loc_sram_buff_w5[164],loc_sram_buff_w5[165],loc_sram_buff_w5[166],loc_sram_buff_w5[167],loc_sram_buff_w5[168],loc_sram_buff_w5[169],loc_sram_buff_w5[170],loc_sram_buff_w5[171],loc_sram_buff_w5[172],loc_sram_buff_w5[173],loc_sram_buff_w5[174],loc_sram_buff_w5[175],loc_sram_buff_w5[176],loc_sram_buff_w5[177],loc_sram_buff_w5[178],loc_sram_buff_w5[179],loc_sram_buff_w5[180],loc_sram_buff_w5[181],loc_sram_buff_w5[182],loc_sram_buff_w5[183],loc_sram_buff_w5[184],loc_sram_buff_w5[185],loc_sram_buff_w5[186],loc_sram_buff_w5[187],loc_sram_buff_w5[188],loc_sram_buff_w5[189],loc_sram_buff_w5[190],loc_sram_buff_w5[191],loc_sram_buff_w5[192],loc_sram_buff_w5[193],loc_sram_buff_w5[194],loc_sram_buff_w5[195],loc_sram_buff_w5[196],loc_sram_buff_w5[197],loc_sram_buff_w5[198],loc_sram_buff_w5[199],loc_sram_buff_w5[200],loc_sram_buff_w5[201],loc_sram_buff_w5[202],loc_sram_buff_w5[203],loc_sram_buff_w5[204],loc_sram_buff_w5[205],loc_sram_buff_w5[206],loc_sram_buff_w5[207],loc_sram_buff_w5[208],loc_sram_buff_w5[209],loc_sram_buff_w5[210],loc_sram_buff_w5[211],loc_sram_buff_w5[212],loc_sram_buff_w5[213],loc_sram_buff_w5[214],loc_sram_buff_w5[215],loc_sram_buff_w5[216],loc_sram_buff_w5[217],loc_sram_buff_w5[218],loc_sram_buff_w5[219],loc_sram_buff_w5[220],loc_sram_buff_w5[221],loc_sram_buff_w5[222],loc_sram_buff_w5[223],loc_sram_buff_w5[224],loc_sram_buff_w5[225],loc_sram_buff_w5[226],loc_sram_buff_w5[227],loc_sram_buff_w5[228],loc_sram_buff_w5[229],loc_sram_buff_w5[230],loc_sram_buff_w5[231],loc_sram_buff_w5[232],loc_sram_buff_w5[233],loc_sram_buff_w5[234],loc_sram_buff_w5[235],loc_sram_buff_w5[236],loc_sram_buff_w5[237],loc_sram_buff_w5[238],loc_sram_buff_w5[239],loc_sram_buff_w5[240],loc_sram_buff_w5[241],loc_sram_buff_w5[242],loc_sram_buff_w5[243],loc_sram_buff_w5[244],loc_sram_buff_w5[245],loc_sram_buff_w5[246],loc_sram_buff_w5[247],loc_sram_buff_w5[248],loc_sram_buff_w5[249],loc_sram_buff_w5[250],loc_sram_buff_w5[251],loc_sram_buff_w5[252],loc_sram_buff_w5[253],loc_sram_buff_w5[254],loc_sram_buff_w5[255]} = loc_sram_rdata5;
	{loc_sram_buff_w6[0],loc_sram_buff_w6[1],loc_sram_buff_w6[2],loc_sram_buff_w6[3],loc_sram_buff_w6[4],loc_sram_buff_w6[5],loc_sram_buff_w6[6],loc_sram_buff_w6[7],loc_sram_buff_w6[8],loc_sram_buff_w6[9],loc_sram_buff_w6[10],loc_sram_buff_w6[11],loc_sram_buff_w6[12],loc_sram_buff_w6[13],loc_sram_buff_w6[14],loc_sram_buff_w6[15],loc_sram_buff_w6[16],loc_sram_buff_w6[17],loc_sram_buff_w6[18],loc_sram_buff_w6[19],loc_sram_buff_w6[20],loc_sram_buff_w6[21],loc_sram_buff_w6[22],loc_sram_buff_w6[23],loc_sram_buff_w6[24],loc_sram_buff_w6[25],loc_sram_buff_w6[26],loc_sram_buff_w6[27],loc_sram_buff_w6[28],loc_sram_buff_w6[29],loc_sram_buff_w6[30],loc_sram_buff_w6[31],loc_sram_buff_w6[32],loc_sram_buff_w6[33],loc_sram_buff_w6[34],loc_sram_buff_w6[35],loc_sram_buff_w6[36],loc_sram_buff_w6[37],loc_sram_buff_w6[38],loc_sram_buff_w6[39],loc_sram_buff_w6[40],loc_sram_buff_w6[41],loc_sram_buff_w6[42],loc_sram_buff_w6[43],loc_sram_buff_w6[44],loc_sram_buff_w6[45],loc_sram_buff_w6[46],loc_sram_buff_w6[47],loc_sram_buff_w6[48],loc_sram_buff_w6[49],loc_sram_buff_w6[50],loc_sram_buff_w6[51],loc_sram_buff_w6[52],loc_sram_buff_w6[53],loc_sram_buff_w6[54],loc_sram_buff_w6[55],loc_sram_buff_w6[56],loc_sram_buff_w6[57],loc_sram_buff_w6[58],loc_sram_buff_w6[59],loc_sram_buff_w6[60],loc_sram_buff_w6[61],loc_sram_buff_w6[62],loc_sram_buff_w6[63],loc_sram_buff_w6[64],loc_sram_buff_w6[65],loc_sram_buff_w6[66],loc_sram_buff_w6[67],loc_sram_buff_w6[68],loc_sram_buff_w6[69],loc_sram_buff_w6[70],loc_sram_buff_w6[71],loc_sram_buff_w6[72],loc_sram_buff_w6[73],loc_sram_buff_w6[74],loc_sram_buff_w6[75],loc_sram_buff_w6[76],loc_sram_buff_w6[77],loc_sram_buff_w6[78],loc_sram_buff_w6[79],loc_sram_buff_w6[80],loc_sram_buff_w6[81],loc_sram_buff_w6[82],loc_sram_buff_w6[83],loc_sram_buff_w6[84],loc_sram_buff_w6[85],loc_sram_buff_w6[86],loc_sram_buff_w6[87],loc_sram_buff_w6[88],loc_sram_buff_w6[89],loc_sram_buff_w6[90],loc_sram_buff_w6[91],loc_sram_buff_w6[92],loc_sram_buff_w6[93],loc_sram_buff_w6[94],loc_sram_buff_w6[95],loc_sram_buff_w6[96],loc_sram_buff_w6[97],loc_sram_buff_w6[98],loc_sram_buff_w6[99],loc_sram_buff_w6[100],loc_sram_buff_w6[101],loc_sram_buff_w6[102],loc_sram_buff_w6[103],loc_sram_buff_w6[104],loc_sram_buff_w6[105],loc_sram_buff_w6[106],loc_sram_buff_w6[107],loc_sram_buff_w6[108],loc_sram_buff_w6[109],loc_sram_buff_w6[110],loc_sram_buff_w6[111],loc_sram_buff_w6[112],loc_sram_buff_w6[113],loc_sram_buff_w6[114],loc_sram_buff_w6[115],loc_sram_buff_w6[116],loc_sram_buff_w6[117],loc_sram_buff_w6[118],loc_sram_buff_w6[119],loc_sram_buff_w6[120],loc_sram_buff_w6[121],loc_sram_buff_w6[122],loc_sram_buff_w6[123],loc_sram_buff_w6[124],loc_sram_buff_w6[125],loc_sram_buff_w6[126],loc_sram_buff_w6[127],loc_sram_buff_w6[128],loc_sram_buff_w6[129],loc_sram_buff_w6[130],loc_sram_buff_w6[131],loc_sram_buff_w6[132],loc_sram_buff_w6[133],loc_sram_buff_w6[134],loc_sram_buff_w6[135],loc_sram_buff_w6[136],loc_sram_buff_w6[137],loc_sram_buff_w6[138],loc_sram_buff_w6[139],loc_sram_buff_w6[140],loc_sram_buff_w6[141],loc_sram_buff_w6[142],loc_sram_buff_w6[143],loc_sram_buff_w6[144],loc_sram_buff_w6[145],loc_sram_buff_w6[146],loc_sram_buff_w6[147],loc_sram_buff_w6[148],loc_sram_buff_w6[149],loc_sram_buff_w6[150],loc_sram_buff_w6[151],loc_sram_buff_w6[152],loc_sram_buff_w6[153],loc_sram_buff_w6[154],loc_sram_buff_w6[155],loc_sram_buff_w6[156],loc_sram_buff_w6[157],loc_sram_buff_w6[158],loc_sram_buff_w6[159],loc_sram_buff_w6[160],loc_sram_buff_w6[161],loc_sram_buff_w6[162],loc_sram_buff_w6[163],loc_sram_buff_w6[164],loc_sram_buff_w6[165],loc_sram_buff_w6[166],loc_sram_buff_w6[167],loc_sram_buff_w6[168],loc_sram_buff_w6[169],loc_sram_buff_w6[170],loc_sram_buff_w6[171],loc_sram_buff_w6[172],loc_sram_buff_w6[173],loc_sram_buff_w6[174],loc_sram_buff_w6[175],loc_sram_buff_w6[176],loc_sram_buff_w6[177],loc_sram_buff_w6[178],loc_sram_buff_w6[179],loc_sram_buff_w6[180],loc_sram_buff_w6[181],loc_sram_buff_w6[182],loc_sram_buff_w6[183],loc_sram_buff_w6[184],loc_sram_buff_w6[185],loc_sram_buff_w6[186],loc_sram_buff_w6[187],loc_sram_buff_w6[188],loc_sram_buff_w6[189],loc_sram_buff_w6[190],loc_sram_buff_w6[191],loc_sram_buff_w6[192],loc_sram_buff_w6[193],loc_sram_buff_w6[194],loc_sram_buff_w6[195],loc_sram_buff_w6[196],loc_sram_buff_w6[197],loc_sram_buff_w6[198],loc_sram_buff_w6[199],loc_sram_buff_w6[200],loc_sram_buff_w6[201],loc_sram_buff_w6[202],loc_sram_buff_w6[203],loc_sram_buff_w6[204],loc_sram_buff_w6[205],loc_sram_buff_w6[206],loc_sram_buff_w6[207],loc_sram_buff_w6[208],loc_sram_buff_w6[209],loc_sram_buff_w6[210],loc_sram_buff_w6[211],loc_sram_buff_w6[212],loc_sram_buff_w6[213],loc_sram_buff_w6[214],loc_sram_buff_w6[215],loc_sram_buff_w6[216],loc_sram_buff_w6[217],loc_sram_buff_w6[218],loc_sram_buff_w6[219],loc_sram_buff_w6[220],loc_sram_buff_w6[221],loc_sram_buff_w6[222],loc_sram_buff_w6[223],loc_sram_buff_w6[224],loc_sram_buff_w6[225],loc_sram_buff_w6[226],loc_sram_buff_w6[227],loc_sram_buff_w6[228],loc_sram_buff_w6[229],loc_sram_buff_w6[230],loc_sram_buff_w6[231],loc_sram_buff_w6[232],loc_sram_buff_w6[233],loc_sram_buff_w6[234],loc_sram_buff_w6[235],loc_sram_buff_w6[236],loc_sram_buff_w6[237],loc_sram_buff_w6[238],loc_sram_buff_w6[239],loc_sram_buff_w6[240],loc_sram_buff_w6[241],loc_sram_buff_w6[242],loc_sram_buff_w6[243],loc_sram_buff_w6[244],loc_sram_buff_w6[245],loc_sram_buff_w6[246],loc_sram_buff_w6[247],loc_sram_buff_w6[248],loc_sram_buff_w6[249],loc_sram_buff_w6[250],loc_sram_buff_w6[251],loc_sram_buff_w6[252],loc_sram_buff_w6[253],loc_sram_buff_w6[254],loc_sram_buff_w6[255]} = loc_sram_rdata6;
	{loc_sram_buff_w7[0],loc_sram_buff_w7[1],loc_sram_buff_w7[2],loc_sram_buff_w7[3],loc_sram_buff_w7[4],loc_sram_buff_w7[5],loc_sram_buff_w7[6],loc_sram_buff_w7[7],loc_sram_buff_w7[8],loc_sram_buff_w7[9],loc_sram_buff_w7[10],loc_sram_buff_w7[11],loc_sram_buff_w7[12],loc_sram_buff_w7[13],loc_sram_buff_w7[14],loc_sram_buff_w7[15],loc_sram_buff_w7[16],loc_sram_buff_w7[17],loc_sram_buff_w7[18],loc_sram_buff_w7[19],loc_sram_buff_w7[20],loc_sram_buff_w7[21],loc_sram_buff_w7[22],loc_sram_buff_w7[23],loc_sram_buff_w7[24],loc_sram_buff_w7[25],loc_sram_buff_w7[26],loc_sram_buff_w7[27],loc_sram_buff_w7[28],loc_sram_buff_w7[29],loc_sram_buff_w7[30],loc_sram_buff_w7[31],loc_sram_buff_w7[32],loc_sram_buff_w7[33],loc_sram_buff_w7[34],loc_sram_buff_w7[35],loc_sram_buff_w7[36],loc_sram_buff_w7[37],loc_sram_buff_w7[38],loc_sram_buff_w7[39],loc_sram_buff_w7[40],loc_sram_buff_w7[41],loc_sram_buff_w7[42],loc_sram_buff_w7[43],loc_sram_buff_w7[44],loc_sram_buff_w7[45],loc_sram_buff_w7[46],loc_sram_buff_w7[47],loc_sram_buff_w7[48],loc_sram_buff_w7[49],loc_sram_buff_w7[50],loc_sram_buff_w7[51],loc_sram_buff_w7[52],loc_sram_buff_w7[53],loc_sram_buff_w7[54],loc_sram_buff_w7[55],loc_sram_buff_w7[56],loc_sram_buff_w7[57],loc_sram_buff_w7[58],loc_sram_buff_w7[59],loc_sram_buff_w7[60],loc_sram_buff_w7[61],loc_sram_buff_w7[62],loc_sram_buff_w7[63],loc_sram_buff_w7[64],loc_sram_buff_w7[65],loc_sram_buff_w7[66],loc_sram_buff_w7[67],loc_sram_buff_w7[68],loc_sram_buff_w7[69],loc_sram_buff_w7[70],loc_sram_buff_w7[71],loc_sram_buff_w7[72],loc_sram_buff_w7[73],loc_sram_buff_w7[74],loc_sram_buff_w7[75],loc_sram_buff_w7[76],loc_sram_buff_w7[77],loc_sram_buff_w7[78],loc_sram_buff_w7[79],loc_sram_buff_w7[80],loc_sram_buff_w7[81],loc_sram_buff_w7[82],loc_sram_buff_w7[83],loc_sram_buff_w7[84],loc_sram_buff_w7[85],loc_sram_buff_w7[86],loc_sram_buff_w7[87],loc_sram_buff_w7[88],loc_sram_buff_w7[89],loc_sram_buff_w7[90],loc_sram_buff_w7[91],loc_sram_buff_w7[92],loc_sram_buff_w7[93],loc_sram_buff_w7[94],loc_sram_buff_w7[95],loc_sram_buff_w7[96],loc_sram_buff_w7[97],loc_sram_buff_w7[98],loc_sram_buff_w7[99],loc_sram_buff_w7[100],loc_sram_buff_w7[101],loc_sram_buff_w7[102],loc_sram_buff_w7[103],loc_sram_buff_w7[104],loc_sram_buff_w7[105],loc_sram_buff_w7[106],loc_sram_buff_w7[107],loc_sram_buff_w7[108],loc_sram_buff_w7[109],loc_sram_buff_w7[110],loc_sram_buff_w7[111],loc_sram_buff_w7[112],loc_sram_buff_w7[113],loc_sram_buff_w7[114],loc_sram_buff_w7[115],loc_sram_buff_w7[116],loc_sram_buff_w7[117],loc_sram_buff_w7[118],loc_sram_buff_w7[119],loc_sram_buff_w7[120],loc_sram_buff_w7[121],loc_sram_buff_w7[122],loc_sram_buff_w7[123],loc_sram_buff_w7[124],loc_sram_buff_w7[125],loc_sram_buff_w7[126],loc_sram_buff_w7[127],loc_sram_buff_w7[128],loc_sram_buff_w7[129],loc_sram_buff_w7[130],loc_sram_buff_w7[131],loc_sram_buff_w7[132],loc_sram_buff_w7[133],loc_sram_buff_w7[134],loc_sram_buff_w7[135],loc_sram_buff_w7[136],loc_sram_buff_w7[137],loc_sram_buff_w7[138],loc_sram_buff_w7[139],loc_sram_buff_w7[140],loc_sram_buff_w7[141],loc_sram_buff_w7[142],loc_sram_buff_w7[143],loc_sram_buff_w7[144],loc_sram_buff_w7[145],loc_sram_buff_w7[146],loc_sram_buff_w7[147],loc_sram_buff_w7[148],loc_sram_buff_w7[149],loc_sram_buff_w7[150],loc_sram_buff_w7[151],loc_sram_buff_w7[152],loc_sram_buff_w7[153],loc_sram_buff_w7[154],loc_sram_buff_w7[155],loc_sram_buff_w7[156],loc_sram_buff_w7[157],loc_sram_buff_w7[158],loc_sram_buff_w7[159],loc_sram_buff_w7[160],loc_sram_buff_w7[161],loc_sram_buff_w7[162],loc_sram_buff_w7[163],loc_sram_buff_w7[164],loc_sram_buff_w7[165],loc_sram_buff_w7[166],loc_sram_buff_w7[167],loc_sram_buff_w7[168],loc_sram_buff_w7[169],loc_sram_buff_w7[170],loc_sram_buff_w7[171],loc_sram_buff_w7[172],loc_sram_buff_w7[173],loc_sram_buff_w7[174],loc_sram_buff_w7[175],loc_sram_buff_w7[176],loc_sram_buff_w7[177],loc_sram_buff_w7[178],loc_sram_buff_w7[179],loc_sram_buff_w7[180],loc_sram_buff_w7[181],loc_sram_buff_w7[182],loc_sram_buff_w7[183],loc_sram_buff_w7[184],loc_sram_buff_w7[185],loc_sram_buff_w7[186],loc_sram_buff_w7[187],loc_sram_buff_w7[188],loc_sram_buff_w7[189],loc_sram_buff_w7[190],loc_sram_buff_w7[191],loc_sram_buff_w7[192],loc_sram_buff_w7[193],loc_sram_buff_w7[194],loc_sram_buff_w7[195],loc_sram_buff_w7[196],loc_sram_buff_w7[197],loc_sram_buff_w7[198],loc_sram_buff_w7[199],loc_sram_buff_w7[200],loc_sram_buff_w7[201],loc_sram_buff_w7[202],loc_sram_buff_w7[203],loc_sram_buff_w7[204],loc_sram_buff_w7[205],loc_sram_buff_w7[206],loc_sram_buff_w7[207],loc_sram_buff_w7[208],loc_sram_buff_w7[209],loc_sram_buff_w7[210],loc_sram_buff_w7[211],loc_sram_buff_w7[212],loc_sram_buff_w7[213],loc_sram_buff_w7[214],loc_sram_buff_w7[215],loc_sram_buff_w7[216],loc_sram_buff_w7[217],loc_sram_buff_w7[218],loc_sram_buff_w7[219],loc_sram_buff_w7[220],loc_sram_buff_w7[221],loc_sram_buff_w7[222],loc_sram_buff_w7[223],loc_sram_buff_w7[224],loc_sram_buff_w7[225],loc_sram_buff_w7[226],loc_sram_buff_w7[227],loc_sram_buff_w7[228],loc_sram_buff_w7[229],loc_sram_buff_w7[230],loc_sram_buff_w7[231],loc_sram_buff_w7[232],loc_sram_buff_w7[233],loc_sram_buff_w7[234],loc_sram_buff_w7[235],loc_sram_buff_w7[236],loc_sram_buff_w7[237],loc_sram_buff_w7[238],loc_sram_buff_w7[239],loc_sram_buff_w7[240],loc_sram_buff_w7[241],loc_sram_buff_w7[242],loc_sram_buff_w7[243],loc_sram_buff_w7[244],loc_sram_buff_w7[245],loc_sram_buff_w7[246],loc_sram_buff_w7[247],loc_sram_buff_w7[248],loc_sram_buff_w7[249],loc_sram_buff_w7[250],loc_sram_buff_w7[251],loc_sram_buff_w7[252],loc_sram_buff_w7[253],loc_sram_buff_w7[254],loc_sram_buff_w7[255]} = loc_sram_rdata7;
	{loc_sram_buff_w8[0],loc_sram_buff_w8[1],loc_sram_buff_w8[2],loc_sram_buff_w8[3],loc_sram_buff_w8[4],loc_sram_buff_w8[5],loc_sram_buff_w8[6],loc_sram_buff_w8[7],loc_sram_buff_w8[8],loc_sram_buff_w8[9],loc_sram_buff_w8[10],loc_sram_buff_w8[11],loc_sram_buff_w8[12],loc_sram_buff_w8[13],loc_sram_buff_w8[14],loc_sram_buff_w8[15],loc_sram_buff_w8[16],loc_sram_buff_w8[17],loc_sram_buff_w8[18],loc_sram_buff_w8[19],loc_sram_buff_w8[20],loc_sram_buff_w8[21],loc_sram_buff_w8[22],loc_sram_buff_w8[23],loc_sram_buff_w8[24],loc_sram_buff_w8[25],loc_sram_buff_w8[26],loc_sram_buff_w8[27],loc_sram_buff_w8[28],loc_sram_buff_w8[29],loc_sram_buff_w8[30],loc_sram_buff_w8[31],loc_sram_buff_w8[32],loc_sram_buff_w8[33],loc_sram_buff_w8[34],loc_sram_buff_w8[35],loc_sram_buff_w8[36],loc_sram_buff_w8[37],loc_sram_buff_w8[38],loc_sram_buff_w8[39],loc_sram_buff_w8[40],loc_sram_buff_w8[41],loc_sram_buff_w8[42],loc_sram_buff_w8[43],loc_sram_buff_w8[44],loc_sram_buff_w8[45],loc_sram_buff_w8[46],loc_sram_buff_w8[47],loc_sram_buff_w8[48],loc_sram_buff_w8[49],loc_sram_buff_w8[50],loc_sram_buff_w8[51],loc_sram_buff_w8[52],loc_sram_buff_w8[53],loc_sram_buff_w8[54],loc_sram_buff_w8[55],loc_sram_buff_w8[56],loc_sram_buff_w8[57],loc_sram_buff_w8[58],loc_sram_buff_w8[59],loc_sram_buff_w8[60],loc_sram_buff_w8[61],loc_sram_buff_w8[62],loc_sram_buff_w8[63],loc_sram_buff_w8[64],loc_sram_buff_w8[65],loc_sram_buff_w8[66],loc_sram_buff_w8[67],loc_sram_buff_w8[68],loc_sram_buff_w8[69],loc_sram_buff_w8[70],loc_sram_buff_w8[71],loc_sram_buff_w8[72],loc_sram_buff_w8[73],loc_sram_buff_w8[74],loc_sram_buff_w8[75],loc_sram_buff_w8[76],loc_sram_buff_w8[77],loc_sram_buff_w8[78],loc_sram_buff_w8[79],loc_sram_buff_w8[80],loc_sram_buff_w8[81],loc_sram_buff_w8[82],loc_sram_buff_w8[83],loc_sram_buff_w8[84],loc_sram_buff_w8[85],loc_sram_buff_w8[86],loc_sram_buff_w8[87],loc_sram_buff_w8[88],loc_sram_buff_w8[89],loc_sram_buff_w8[90],loc_sram_buff_w8[91],loc_sram_buff_w8[92],loc_sram_buff_w8[93],loc_sram_buff_w8[94],loc_sram_buff_w8[95],loc_sram_buff_w8[96],loc_sram_buff_w8[97],loc_sram_buff_w8[98],loc_sram_buff_w8[99],loc_sram_buff_w8[100],loc_sram_buff_w8[101],loc_sram_buff_w8[102],loc_sram_buff_w8[103],loc_sram_buff_w8[104],loc_sram_buff_w8[105],loc_sram_buff_w8[106],loc_sram_buff_w8[107],loc_sram_buff_w8[108],loc_sram_buff_w8[109],loc_sram_buff_w8[110],loc_sram_buff_w8[111],loc_sram_buff_w8[112],loc_sram_buff_w8[113],loc_sram_buff_w8[114],loc_sram_buff_w8[115],loc_sram_buff_w8[116],loc_sram_buff_w8[117],loc_sram_buff_w8[118],loc_sram_buff_w8[119],loc_sram_buff_w8[120],loc_sram_buff_w8[121],loc_sram_buff_w8[122],loc_sram_buff_w8[123],loc_sram_buff_w8[124],loc_sram_buff_w8[125],loc_sram_buff_w8[126],loc_sram_buff_w8[127],loc_sram_buff_w8[128],loc_sram_buff_w8[129],loc_sram_buff_w8[130],loc_sram_buff_w8[131],loc_sram_buff_w8[132],loc_sram_buff_w8[133],loc_sram_buff_w8[134],loc_sram_buff_w8[135],loc_sram_buff_w8[136],loc_sram_buff_w8[137],loc_sram_buff_w8[138],loc_sram_buff_w8[139],loc_sram_buff_w8[140],loc_sram_buff_w8[141],loc_sram_buff_w8[142],loc_sram_buff_w8[143],loc_sram_buff_w8[144],loc_sram_buff_w8[145],loc_sram_buff_w8[146],loc_sram_buff_w8[147],loc_sram_buff_w8[148],loc_sram_buff_w8[149],loc_sram_buff_w8[150],loc_sram_buff_w8[151],loc_sram_buff_w8[152],loc_sram_buff_w8[153],loc_sram_buff_w8[154],loc_sram_buff_w8[155],loc_sram_buff_w8[156],loc_sram_buff_w8[157],loc_sram_buff_w8[158],loc_sram_buff_w8[159],loc_sram_buff_w8[160],loc_sram_buff_w8[161],loc_sram_buff_w8[162],loc_sram_buff_w8[163],loc_sram_buff_w8[164],loc_sram_buff_w8[165],loc_sram_buff_w8[166],loc_sram_buff_w8[167],loc_sram_buff_w8[168],loc_sram_buff_w8[169],loc_sram_buff_w8[170],loc_sram_buff_w8[171],loc_sram_buff_w8[172],loc_sram_buff_w8[173],loc_sram_buff_w8[174],loc_sram_buff_w8[175],loc_sram_buff_w8[176],loc_sram_buff_w8[177],loc_sram_buff_w8[178],loc_sram_buff_w8[179],loc_sram_buff_w8[180],loc_sram_buff_w8[181],loc_sram_buff_w8[182],loc_sram_buff_w8[183],loc_sram_buff_w8[184],loc_sram_buff_w8[185],loc_sram_buff_w8[186],loc_sram_buff_w8[187],loc_sram_buff_w8[188],loc_sram_buff_w8[189],loc_sram_buff_w8[190],loc_sram_buff_w8[191],loc_sram_buff_w8[192],loc_sram_buff_w8[193],loc_sram_buff_w8[194],loc_sram_buff_w8[195],loc_sram_buff_w8[196],loc_sram_buff_w8[197],loc_sram_buff_w8[198],loc_sram_buff_w8[199],loc_sram_buff_w8[200],loc_sram_buff_w8[201],loc_sram_buff_w8[202],loc_sram_buff_w8[203],loc_sram_buff_w8[204],loc_sram_buff_w8[205],loc_sram_buff_w8[206],loc_sram_buff_w8[207],loc_sram_buff_w8[208],loc_sram_buff_w8[209],loc_sram_buff_w8[210],loc_sram_buff_w8[211],loc_sram_buff_w8[212],loc_sram_buff_w8[213],loc_sram_buff_w8[214],loc_sram_buff_w8[215],loc_sram_buff_w8[216],loc_sram_buff_w8[217],loc_sram_buff_w8[218],loc_sram_buff_w8[219],loc_sram_buff_w8[220],loc_sram_buff_w8[221],loc_sram_buff_w8[222],loc_sram_buff_w8[223],loc_sram_buff_w8[224],loc_sram_buff_w8[225],loc_sram_buff_w8[226],loc_sram_buff_w8[227],loc_sram_buff_w8[228],loc_sram_buff_w8[229],loc_sram_buff_w8[230],loc_sram_buff_w8[231],loc_sram_buff_w8[232],loc_sram_buff_w8[233],loc_sram_buff_w8[234],loc_sram_buff_w8[235],loc_sram_buff_w8[236],loc_sram_buff_w8[237],loc_sram_buff_w8[238],loc_sram_buff_w8[239],loc_sram_buff_w8[240],loc_sram_buff_w8[241],loc_sram_buff_w8[242],loc_sram_buff_w8[243],loc_sram_buff_w8[244],loc_sram_buff_w8[245],loc_sram_buff_w8[246],loc_sram_buff_w8[247],loc_sram_buff_w8[248],loc_sram_buff_w8[249],loc_sram_buff_w8[250],loc_sram_buff_w8[251],loc_sram_buff_w8[252],loc_sram_buff_w8[253],loc_sram_buff_w8[254],loc_sram_buff_w8[255]} = loc_sram_rdata8;
	{loc_sram_buff_w9[0],loc_sram_buff_w9[1],loc_sram_buff_w9[2],loc_sram_buff_w9[3],loc_sram_buff_w9[4],loc_sram_buff_w9[5],loc_sram_buff_w9[6],loc_sram_buff_w9[7],loc_sram_buff_w9[8],loc_sram_buff_w9[9],loc_sram_buff_w9[10],loc_sram_buff_w9[11],loc_sram_buff_w9[12],loc_sram_buff_w9[13],loc_sram_buff_w9[14],loc_sram_buff_w9[15],loc_sram_buff_w9[16],loc_sram_buff_w9[17],loc_sram_buff_w9[18],loc_sram_buff_w9[19],loc_sram_buff_w9[20],loc_sram_buff_w9[21],loc_sram_buff_w9[22],loc_sram_buff_w9[23],loc_sram_buff_w9[24],loc_sram_buff_w9[25],loc_sram_buff_w9[26],loc_sram_buff_w9[27],loc_sram_buff_w9[28],loc_sram_buff_w9[29],loc_sram_buff_w9[30],loc_sram_buff_w9[31],loc_sram_buff_w9[32],loc_sram_buff_w9[33],loc_sram_buff_w9[34],loc_sram_buff_w9[35],loc_sram_buff_w9[36],loc_sram_buff_w9[37],loc_sram_buff_w9[38],loc_sram_buff_w9[39],loc_sram_buff_w9[40],loc_sram_buff_w9[41],loc_sram_buff_w9[42],loc_sram_buff_w9[43],loc_sram_buff_w9[44],loc_sram_buff_w9[45],loc_sram_buff_w9[46],loc_sram_buff_w9[47],loc_sram_buff_w9[48],loc_sram_buff_w9[49],loc_sram_buff_w9[50],loc_sram_buff_w9[51],loc_sram_buff_w9[52],loc_sram_buff_w9[53],loc_sram_buff_w9[54],loc_sram_buff_w9[55],loc_sram_buff_w9[56],loc_sram_buff_w9[57],loc_sram_buff_w9[58],loc_sram_buff_w9[59],loc_sram_buff_w9[60],loc_sram_buff_w9[61],loc_sram_buff_w9[62],loc_sram_buff_w9[63],loc_sram_buff_w9[64],loc_sram_buff_w9[65],loc_sram_buff_w9[66],loc_sram_buff_w9[67],loc_sram_buff_w9[68],loc_sram_buff_w9[69],loc_sram_buff_w9[70],loc_sram_buff_w9[71],loc_sram_buff_w9[72],loc_sram_buff_w9[73],loc_sram_buff_w9[74],loc_sram_buff_w9[75],loc_sram_buff_w9[76],loc_sram_buff_w9[77],loc_sram_buff_w9[78],loc_sram_buff_w9[79],loc_sram_buff_w9[80],loc_sram_buff_w9[81],loc_sram_buff_w9[82],loc_sram_buff_w9[83],loc_sram_buff_w9[84],loc_sram_buff_w9[85],loc_sram_buff_w9[86],loc_sram_buff_w9[87],loc_sram_buff_w9[88],loc_sram_buff_w9[89],loc_sram_buff_w9[90],loc_sram_buff_w9[91],loc_sram_buff_w9[92],loc_sram_buff_w9[93],loc_sram_buff_w9[94],loc_sram_buff_w9[95],loc_sram_buff_w9[96],loc_sram_buff_w9[97],loc_sram_buff_w9[98],loc_sram_buff_w9[99],loc_sram_buff_w9[100],loc_sram_buff_w9[101],loc_sram_buff_w9[102],loc_sram_buff_w9[103],loc_sram_buff_w9[104],loc_sram_buff_w9[105],loc_sram_buff_w9[106],loc_sram_buff_w9[107],loc_sram_buff_w9[108],loc_sram_buff_w9[109],loc_sram_buff_w9[110],loc_sram_buff_w9[111],loc_sram_buff_w9[112],loc_sram_buff_w9[113],loc_sram_buff_w9[114],loc_sram_buff_w9[115],loc_sram_buff_w9[116],loc_sram_buff_w9[117],loc_sram_buff_w9[118],loc_sram_buff_w9[119],loc_sram_buff_w9[120],loc_sram_buff_w9[121],loc_sram_buff_w9[122],loc_sram_buff_w9[123],loc_sram_buff_w9[124],loc_sram_buff_w9[125],loc_sram_buff_w9[126],loc_sram_buff_w9[127],loc_sram_buff_w9[128],loc_sram_buff_w9[129],loc_sram_buff_w9[130],loc_sram_buff_w9[131],loc_sram_buff_w9[132],loc_sram_buff_w9[133],loc_sram_buff_w9[134],loc_sram_buff_w9[135],loc_sram_buff_w9[136],loc_sram_buff_w9[137],loc_sram_buff_w9[138],loc_sram_buff_w9[139],loc_sram_buff_w9[140],loc_sram_buff_w9[141],loc_sram_buff_w9[142],loc_sram_buff_w9[143],loc_sram_buff_w9[144],loc_sram_buff_w9[145],loc_sram_buff_w9[146],loc_sram_buff_w9[147],loc_sram_buff_w9[148],loc_sram_buff_w9[149],loc_sram_buff_w9[150],loc_sram_buff_w9[151],loc_sram_buff_w9[152],loc_sram_buff_w9[153],loc_sram_buff_w9[154],loc_sram_buff_w9[155],loc_sram_buff_w9[156],loc_sram_buff_w9[157],loc_sram_buff_w9[158],loc_sram_buff_w9[159],loc_sram_buff_w9[160],loc_sram_buff_w9[161],loc_sram_buff_w9[162],loc_sram_buff_w9[163],loc_sram_buff_w9[164],loc_sram_buff_w9[165],loc_sram_buff_w9[166],loc_sram_buff_w9[167],loc_sram_buff_w9[168],loc_sram_buff_w9[169],loc_sram_buff_w9[170],loc_sram_buff_w9[171],loc_sram_buff_w9[172],loc_sram_buff_w9[173],loc_sram_buff_w9[174],loc_sram_buff_w9[175],loc_sram_buff_w9[176],loc_sram_buff_w9[177],loc_sram_buff_w9[178],loc_sram_buff_w9[179],loc_sram_buff_w9[180],loc_sram_buff_w9[181],loc_sram_buff_w9[182],loc_sram_buff_w9[183],loc_sram_buff_w9[184],loc_sram_buff_w9[185],loc_sram_buff_w9[186],loc_sram_buff_w9[187],loc_sram_buff_w9[188],loc_sram_buff_w9[189],loc_sram_buff_w9[190],loc_sram_buff_w9[191],loc_sram_buff_w9[192],loc_sram_buff_w9[193],loc_sram_buff_w9[194],loc_sram_buff_w9[195],loc_sram_buff_w9[196],loc_sram_buff_w9[197],loc_sram_buff_w9[198],loc_sram_buff_w9[199],loc_sram_buff_w9[200],loc_sram_buff_w9[201],loc_sram_buff_w9[202],loc_sram_buff_w9[203],loc_sram_buff_w9[204],loc_sram_buff_w9[205],loc_sram_buff_w9[206],loc_sram_buff_w9[207],loc_sram_buff_w9[208],loc_sram_buff_w9[209],loc_sram_buff_w9[210],loc_sram_buff_w9[211],loc_sram_buff_w9[212],loc_sram_buff_w9[213],loc_sram_buff_w9[214],loc_sram_buff_w9[215],loc_sram_buff_w9[216],loc_sram_buff_w9[217],loc_sram_buff_w9[218],loc_sram_buff_w9[219],loc_sram_buff_w9[220],loc_sram_buff_w9[221],loc_sram_buff_w9[222],loc_sram_buff_w9[223],loc_sram_buff_w9[224],loc_sram_buff_w9[225],loc_sram_buff_w9[226],loc_sram_buff_w9[227],loc_sram_buff_w9[228],loc_sram_buff_w9[229],loc_sram_buff_w9[230],loc_sram_buff_w9[231],loc_sram_buff_w9[232],loc_sram_buff_w9[233],loc_sram_buff_w9[234],loc_sram_buff_w9[235],loc_sram_buff_w9[236],loc_sram_buff_w9[237],loc_sram_buff_w9[238],loc_sram_buff_w9[239],loc_sram_buff_w9[240],loc_sram_buff_w9[241],loc_sram_buff_w9[242],loc_sram_buff_w9[243],loc_sram_buff_w9[244],loc_sram_buff_w9[245],loc_sram_buff_w9[246],loc_sram_buff_w9[247],loc_sram_buff_w9[248],loc_sram_buff_w9[249],loc_sram_buff_w9[250],loc_sram_buff_w9[251],loc_sram_buff_w9[252],loc_sram_buff_w9[253],loc_sram_buff_w9[254],loc_sram_buff_w9[255]} = loc_sram_rdata9;
	{loc_sram_buff_w10[0],loc_sram_buff_w10[1],loc_sram_buff_w10[2],loc_sram_buff_w10[3],loc_sram_buff_w10[4],loc_sram_buff_w10[5],loc_sram_buff_w10[6],loc_sram_buff_w10[7],loc_sram_buff_w10[8],loc_sram_buff_w10[9],loc_sram_buff_w10[10],loc_sram_buff_w10[11],loc_sram_buff_w10[12],loc_sram_buff_w10[13],loc_sram_buff_w10[14],loc_sram_buff_w10[15],loc_sram_buff_w10[16],loc_sram_buff_w10[17],loc_sram_buff_w10[18],loc_sram_buff_w10[19],loc_sram_buff_w10[20],loc_sram_buff_w10[21],loc_sram_buff_w10[22],loc_sram_buff_w10[23],loc_sram_buff_w10[24],loc_sram_buff_w10[25],loc_sram_buff_w10[26],loc_sram_buff_w10[27],loc_sram_buff_w10[28],loc_sram_buff_w10[29],loc_sram_buff_w10[30],loc_sram_buff_w10[31],loc_sram_buff_w10[32],loc_sram_buff_w10[33],loc_sram_buff_w10[34],loc_sram_buff_w10[35],loc_sram_buff_w10[36],loc_sram_buff_w10[37],loc_sram_buff_w10[38],loc_sram_buff_w10[39],loc_sram_buff_w10[40],loc_sram_buff_w10[41],loc_sram_buff_w10[42],loc_sram_buff_w10[43],loc_sram_buff_w10[44],loc_sram_buff_w10[45],loc_sram_buff_w10[46],loc_sram_buff_w10[47],loc_sram_buff_w10[48],loc_sram_buff_w10[49],loc_sram_buff_w10[50],loc_sram_buff_w10[51],loc_sram_buff_w10[52],loc_sram_buff_w10[53],loc_sram_buff_w10[54],loc_sram_buff_w10[55],loc_sram_buff_w10[56],loc_sram_buff_w10[57],loc_sram_buff_w10[58],loc_sram_buff_w10[59],loc_sram_buff_w10[60],loc_sram_buff_w10[61],loc_sram_buff_w10[62],loc_sram_buff_w10[63],loc_sram_buff_w10[64],loc_sram_buff_w10[65],loc_sram_buff_w10[66],loc_sram_buff_w10[67],loc_sram_buff_w10[68],loc_sram_buff_w10[69],loc_sram_buff_w10[70],loc_sram_buff_w10[71],loc_sram_buff_w10[72],loc_sram_buff_w10[73],loc_sram_buff_w10[74],loc_sram_buff_w10[75],loc_sram_buff_w10[76],loc_sram_buff_w10[77],loc_sram_buff_w10[78],loc_sram_buff_w10[79],loc_sram_buff_w10[80],loc_sram_buff_w10[81],loc_sram_buff_w10[82],loc_sram_buff_w10[83],loc_sram_buff_w10[84],loc_sram_buff_w10[85],loc_sram_buff_w10[86],loc_sram_buff_w10[87],loc_sram_buff_w10[88],loc_sram_buff_w10[89],loc_sram_buff_w10[90],loc_sram_buff_w10[91],loc_sram_buff_w10[92],loc_sram_buff_w10[93],loc_sram_buff_w10[94],loc_sram_buff_w10[95],loc_sram_buff_w10[96],loc_sram_buff_w10[97],loc_sram_buff_w10[98],loc_sram_buff_w10[99],loc_sram_buff_w10[100],loc_sram_buff_w10[101],loc_sram_buff_w10[102],loc_sram_buff_w10[103],loc_sram_buff_w10[104],loc_sram_buff_w10[105],loc_sram_buff_w10[106],loc_sram_buff_w10[107],loc_sram_buff_w10[108],loc_sram_buff_w10[109],loc_sram_buff_w10[110],loc_sram_buff_w10[111],loc_sram_buff_w10[112],loc_sram_buff_w10[113],loc_sram_buff_w10[114],loc_sram_buff_w10[115],loc_sram_buff_w10[116],loc_sram_buff_w10[117],loc_sram_buff_w10[118],loc_sram_buff_w10[119],loc_sram_buff_w10[120],loc_sram_buff_w10[121],loc_sram_buff_w10[122],loc_sram_buff_w10[123],loc_sram_buff_w10[124],loc_sram_buff_w10[125],loc_sram_buff_w10[126],loc_sram_buff_w10[127],loc_sram_buff_w10[128],loc_sram_buff_w10[129],loc_sram_buff_w10[130],loc_sram_buff_w10[131],loc_sram_buff_w10[132],loc_sram_buff_w10[133],loc_sram_buff_w10[134],loc_sram_buff_w10[135],loc_sram_buff_w10[136],loc_sram_buff_w10[137],loc_sram_buff_w10[138],loc_sram_buff_w10[139],loc_sram_buff_w10[140],loc_sram_buff_w10[141],loc_sram_buff_w10[142],loc_sram_buff_w10[143],loc_sram_buff_w10[144],loc_sram_buff_w10[145],loc_sram_buff_w10[146],loc_sram_buff_w10[147],loc_sram_buff_w10[148],loc_sram_buff_w10[149],loc_sram_buff_w10[150],loc_sram_buff_w10[151],loc_sram_buff_w10[152],loc_sram_buff_w10[153],loc_sram_buff_w10[154],loc_sram_buff_w10[155],loc_sram_buff_w10[156],loc_sram_buff_w10[157],loc_sram_buff_w10[158],loc_sram_buff_w10[159],loc_sram_buff_w10[160],loc_sram_buff_w10[161],loc_sram_buff_w10[162],loc_sram_buff_w10[163],loc_sram_buff_w10[164],loc_sram_buff_w10[165],loc_sram_buff_w10[166],loc_sram_buff_w10[167],loc_sram_buff_w10[168],loc_sram_buff_w10[169],loc_sram_buff_w10[170],loc_sram_buff_w10[171],loc_sram_buff_w10[172],loc_sram_buff_w10[173],loc_sram_buff_w10[174],loc_sram_buff_w10[175],loc_sram_buff_w10[176],loc_sram_buff_w10[177],loc_sram_buff_w10[178],loc_sram_buff_w10[179],loc_sram_buff_w10[180],loc_sram_buff_w10[181],loc_sram_buff_w10[182],loc_sram_buff_w10[183],loc_sram_buff_w10[184],loc_sram_buff_w10[185],loc_sram_buff_w10[186],loc_sram_buff_w10[187],loc_sram_buff_w10[188],loc_sram_buff_w10[189],loc_sram_buff_w10[190],loc_sram_buff_w10[191],loc_sram_buff_w10[192],loc_sram_buff_w10[193],loc_sram_buff_w10[194],loc_sram_buff_w10[195],loc_sram_buff_w10[196],loc_sram_buff_w10[197],loc_sram_buff_w10[198],loc_sram_buff_w10[199],loc_sram_buff_w10[200],loc_sram_buff_w10[201],loc_sram_buff_w10[202],loc_sram_buff_w10[203],loc_sram_buff_w10[204],loc_sram_buff_w10[205],loc_sram_buff_w10[206],loc_sram_buff_w10[207],loc_sram_buff_w10[208],loc_sram_buff_w10[209],loc_sram_buff_w10[210],loc_sram_buff_w10[211],loc_sram_buff_w10[212],loc_sram_buff_w10[213],loc_sram_buff_w10[214],loc_sram_buff_w10[215],loc_sram_buff_w10[216],loc_sram_buff_w10[217],loc_sram_buff_w10[218],loc_sram_buff_w10[219],loc_sram_buff_w10[220],loc_sram_buff_w10[221],loc_sram_buff_w10[222],loc_sram_buff_w10[223],loc_sram_buff_w10[224],loc_sram_buff_w10[225],loc_sram_buff_w10[226],loc_sram_buff_w10[227],loc_sram_buff_w10[228],loc_sram_buff_w10[229],loc_sram_buff_w10[230],loc_sram_buff_w10[231],loc_sram_buff_w10[232],loc_sram_buff_w10[233],loc_sram_buff_w10[234],loc_sram_buff_w10[235],loc_sram_buff_w10[236],loc_sram_buff_w10[237],loc_sram_buff_w10[238],loc_sram_buff_w10[239],loc_sram_buff_w10[240],loc_sram_buff_w10[241],loc_sram_buff_w10[242],loc_sram_buff_w10[243],loc_sram_buff_w10[244],loc_sram_buff_w10[245],loc_sram_buff_w10[246],loc_sram_buff_w10[247],loc_sram_buff_w10[248],loc_sram_buff_w10[249],loc_sram_buff_w10[250],loc_sram_buff_w10[251],loc_sram_buff_w10[252],loc_sram_buff_w10[253],loc_sram_buff_w10[254],loc_sram_buff_w10[255]} = loc_sram_rdata10;
	{loc_sram_buff_w11[0],loc_sram_buff_w11[1],loc_sram_buff_w11[2],loc_sram_buff_w11[3],loc_sram_buff_w11[4],loc_sram_buff_w11[5],loc_sram_buff_w11[6],loc_sram_buff_w11[7],loc_sram_buff_w11[8],loc_sram_buff_w11[9],loc_sram_buff_w11[10],loc_sram_buff_w11[11],loc_sram_buff_w11[12],loc_sram_buff_w11[13],loc_sram_buff_w11[14],loc_sram_buff_w11[15],loc_sram_buff_w11[16],loc_sram_buff_w11[17],loc_sram_buff_w11[18],loc_sram_buff_w11[19],loc_sram_buff_w11[20],loc_sram_buff_w11[21],loc_sram_buff_w11[22],loc_sram_buff_w11[23],loc_sram_buff_w11[24],loc_sram_buff_w11[25],loc_sram_buff_w11[26],loc_sram_buff_w11[27],loc_sram_buff_w11[28],loc_sram_buff_w11[29],loc_sram_buff_w11[30],loc_sram_buff_w11[31],loc_sram_buff_w11[32],loc_sram_buff_w11[33],loc_sram_buff_w11[34],loc_sram_buff_w11[35],loc_sram_buff_w11[36],loc_sram_buff_w11[37],loc_sram_buff_w11[38],loc_sram_buff_w11[39],loc_sram_buff_w11[40],loc_sram_buff_w11[41],loc_sram_buff_w11[42],loc_sram_buff_w11[43],loc_sram_buff_w11[44],loc_sram_buff_w11[45],loc_sram_buff_w11[46],loc_sram_buff_w11[47],loc_sram_buff_w11[48],loc_sram_buff_w11[49],loc_sram_buff_w11[50],loc_sram_buff_w11[51],loc_sram_buff_w11[52],loc_sram_buff_w11[53],loc_sram_buff_w11[54],loc_sram_buff_w11[55],loc_sram_buff_w11[56],loc_sram_buff_w11[57],loc_sram_buff_w11[58],loc_sram_buff_w11[59],loc_sram_buff_w11[60],loc_sram_buff_w11[61],loc_sram_buff_w11[62],loc_sram_buff_w11[63],loc_sram_buff_w11[64],loc_sram_buff_w11[65],loc_sram_buff_w11[66],loc_sram_buff_w11[67],loc_sram_buff_w11[68],loc_sram_buff_w11[69],loc_sram_buff_w11[70],loc_sram_buff_w11[71],loc_sram_buff_w11[72],loc_sram_buff_w11[73],loc_sram_buff_w11[74],loc_sram_buff_w11[75],loc_sram_buff_w11[76],loc_sram_buff_w11[77],loc_sram_buff_w11[78],loc_sram_buff_w11[79],loc_sram_buff_w11[80],loc_sram_buff_w11[81],loc_sram_buff_w11[82],loc_sram_buff_w11[83],loc_sram_buff_w11[84],loc_sram_buff_w11[85],loc_sram_buff_w11[86],loc_sram_buff_w11[87],loc_sram_buff_w11[88],loc_sram_buff_w11[89],loc_sram_buff_w11[90],loc_sram_buff_w11[91],loc_sram_buff_w11[92],loc_sram_buff_w11[93],loc_sram_buff_w11[94],loc_sram_buff_w11[95],loc_sram_buff_w11[96],loc_sram_buff_w11[97],loc_sram_buff_w11[98],loc_sram_buff_w11[99],loc_sram_buff_w11[100],loc_sram_buff_w11[101],loc_sram_buff_w11[102],loc_sram_buff_w11[103],loc_sram_buff_w11[104],loc_sram_buff_w11[105],loc_sram_buff_w11[106],loc_sram_buff_w11[107],loc_sram_buff_w11[108],loc_sram_buff_w11[109],loc_sram_buff_w11[110],loc_sram_buff_w11[111],loc_sram_buff_w11[112],loc_sram_buff_w11[113],loc_sram_buff_w11[114],loc_sram_buff_w11[115],loc_sram_buff_w11[116],loc_sram_buff_w11[117],loc_sram_buff_w11[118],loc_sram_buff_w11[119],loc_sram_buff_w11[120],loc_sram_buff_w11[121],loc_sram_buff_w11[122],loc_sram_buff_w11[123],loc_sram_buff_w11[124],loc_sram_buff_w11[125],loc_sram_buff_w11[126],loc_sram_buff_w11[127],loc_sram_buff_w11[128],loc_sram_buff_w11[129],loc_sram_buff_w11[130],loc_sram_buff_w11[131],loc_sram_buff_w11[132],loc_sram_buff_w11[133],loc_sram_buff_w11[134],loc_sram_buff_w11[135],loc_sram_buff_w11[136],loc_sram_buff_w11[137],loc_sram_buff_w11[138],loc_sram_buff_w11[139],loc_sram_buff_w11[140],loc_sram_buff_w11[141],loc_sram_buff_w11[142],loc_sram_buff_w11[143],loc_sram_buff_w11[144],loc_sram_buff_w11[145],loc_sram_buff_w11[146],loc_sram_buff_w11[147],loc_sram_buff_w11[148],loc_sram_buff_w11[149],loc_sram_buff_w11[150],loc_sram_buff_w11[151],loc_sram_buff_w11[152],loc_sram_buff_w11[153],loc_sram_buff_w11[154],loc_sram_buff_w11[155],loc_sram_buff_w11[156],loc_sram_buff_w11[157],loc_sram_buff_w11[158],loc_sram_buff_w11[159],loc_sram_buff_w11[160],loc_sram_buff_w11[161],loc_sram_buff_w11[162],loc_sram_buff_w11[163],loc_sram_buff_w11[164],loc_sram_buff_w11[165],loc_sram_buff_w11[166],loc_sram_buff_w11[167],loc_sram_buff_w11[168],loc_sram_buff_w11[169],loc_sram_buff_w11[170],loc_sram_buff_w11[171],loc_sram_buff_w11[172],loc_sram_buff_w11[173],loc_sram_buff_w11[174],loc_sram_buff_w11[175],loc_sram_buff_w11[176],loc_sram_buff_w11[177],loc_sram_buff_w11[178],loc_sram_buff_w11[179],loc_sram_buff_w11[180],loc_sram_buff_w11[181],loc_sram_buff_w11[182],loc_sram_buff_w11[183],loc_sram_buff_w11[184],loc_sram_buff_w11[185],loc_sram_buff_w11[186],loc_sram_buff_w11[187],loc_sram_buff_w11[188],loc_sram_buff_w11[189],loc_sram_buff_w11[190],loc_sram_buff_w11[191],loc_sram_buff_w11[192],loc_sram_buff_w11[193],loc_sram_buff_w11[194],loc_sram_buff_w11[195],loc_sram_buff_w11[196],loc_sram_buff_w11[197],loc_sram_buff_w11[198],loc_sram_buff_w11[199],loc_sram_buff_w11[200],loc_sram_buff_w11[201],loc_sram_buff_w11[202],loc_sram_buff_w11[203],loc_sram_buff_w11[204],loc_sram_buff_w11[205],loc_sram_buff_w11[206],loc_sram_buff_w11[207],loc_sram_buff_w11[208],loc_sram_buff_w11[209],loc_sram_buff_w11[210],loc_sram_buff_w11[211],loc_sram_buff_w11[212],loc_sram_buff_w11[213],loc_sram_buff_w11[214],loc_sram_buff_w11[215],loc_sram_buff_w11[216],loc_sram_buff_w11[217],loc_sram_buff_w11[218],loc_sram_buff_w11[219],loc_sram_buff_w11[220],loc_sram_buff_w11[221],loc_sram_buff_w11[222],loc_sram_buff_w11[223],loc_sram_buff_w11[224],loc_sram_buff_w11[225],loc_sram_buff_w11[226],loc_sram_buff_w11[227],loc_sram_buff_w11[228],loc_sram_buff_w11[229],loc_sram_buff_w11[230],loc_sram_buff_w11[231],loc_sram_buff_w11[232],loc_sram_buff_w11[233],loc_sram_buff_w11[234],loc_sram_buff_w11[235],loc_sram_buff_w11[236],loc_sram_buff_w11[237],loc_sram_buff_w11[238],loc_sram_buff_w11[239],loc_sram_buff_w11[240],loc_sram_buff_w11[241],loc_sram_buff_w11[242],loc_sram_buff_w11[243],loc_sram_buff_w11[244],loc_sram_buff_w11[245],loc_sram_buff_w11[246],loc_sram_buff_w11[247],loc_sram_buff_w11[248],loc_sram_buff_w11[249],loc_sram_buff_w11[250],loc_sram_buff_w11[251],loc_sram_buff_w11[252],loc_sram_buff_w11[253],loc_sram_buff_w11[254],loc_sram_buff_w11[255]} = loc_sram_rdata11;
	{loc_sram_buff_w12[0],loc_sram_buff_w12[1],loc_sram_buff_w12[2],loc_sram_buff_w12[3],loc_sram_buff_w12[4],loc_sram_buff_w12[5],loc_sram_buff_w12[6],loc_sram_buff_w12[7],loc_sram_buff_w12[8],loc_sram_buff_w12[9],loc_sram_buff_w12[10],loc_sram_buff_w12[11],loc_sram_buff_w12[12],loc_sram_buff_w12[13],loc_sram_buff_w12[14],loc_sram_buff_w12[15],loc_sram_buff_w12[16],loc_sram_buff_w12[17],loc_sram_buff_w12[18],loc_sram_buff_w12[19],loc_sram_buff_w12[20],loc_sram_buff_w12[21],loc_sram_buff_w12[22],loc_sram_buff_w12[23],loc_sram_buff_w12[24],loc_sram_buff_w12[25],loc_sram_buff_w12[26],loc_sram_buff_w12[27],loc_sram_buff_w12[28],loc_sram_buff_w12[29],loc_sram_buff_w12[30],loc_sram_buff_w12[31],loc_sram_buff_w12[32],loc_sram_buff_w12[33],loc_sram_buff_w12[34],loc_sram_buff_w12[35],loc_sram_buff_w12[36],loc_sram_buff_w12[37],loc_sram_buff_w12[38],loc_sram_buff_w12[39],loc_sram_buff_w12[40],loc_sram_buff_w12[41],loc_sram_buff_w12[42],loc_sram_buff_w12[43],loc_sram_buff_w12[44],loc_sram_buff_w12[45],loc_sram_buff_w12[46],loc_sram_buff_w12[47],loc_sram_buff_w12[48],loc_sram_buff_w12[49],loc_sram_buff_w12[50],loc_sram_buff_w12[51],loc_sram_buff_w12[52],loc_sram_buff_w12[53],loc_sram_buff_w12[54],loc_sram_buff_w12[55],loc_sram_buff_w12[56],loc_sram_buff_w12[57],loc_sram_buff_w12[58],loc_sram_buff_w12[59],loc_sram_buff_w12[60],loc_sram_buff_w12[61],loc_sram_buff_w12[62],loc_sram_buff_w12[63],loc_sram_buff_w12[64],loc_sram_buff_w12[65],loc_sram_buff_w12[66],loc_sram_buff_w12[67],loc_sram_buff_w12[68],loc_sram_buff_w12[69],loc_sram_buff_w12[70],loc_sram_buff_w12[71],loc_sram_buff_w12[72],loc_sram_buff_w12[73],loc_sram_buff_w12[74],loc_sram_buff_w12[75],loc_sram_buff_w12[76],loc_sram_buff_w12[77],loc_sram_buff_w12[78],loc_sram_buff_w12[79],loc_sram_buff_w12[80],loc_sram_buff_w12[81],loc_sram_buff_w12[82],loc_sram_buff_w12[83],loc_sram_buff_w12[84],loc_sram_buff_w12[85],loc_sram_buff_w12[86],loc_sram_buff_w12[87],loc_sram_buff_w12[88],loc_sram_buff_w12[89],loc_sram_buff_w12[90],loc_sram_buff_w12[91],loc_sram_buff_w12[92],loc_sram_buff_w12[93],loc_sram_buff_w12[94],loc_sram_buff_w12[95],loc_sram_buff_w12[96],loc_sram_buff_w12[97],loc_sram_buff_w12[98],loc_sram_buff_w12[99],loc_sram_buff_w12[100],loc_sram_buff_w12[101],loc_sram_buff_w12[102],loc_sram_buff_w12[103],loc_sram_buff_w12[104],loc_sram_buff_w12[105],loc_sram_buff_w12[106],loc_sram_buff_w12[107],loc_sram_buff_w12[108],loc_sram_buff_w12[109],loc_sram_buff_w12[110],loc_sram_buff_w12[111],loc_sram_buff_w12[112],loc_sram_buff_w12[113],loc_sram_buff_w12[114],loc_sram_buff_w12[115],loc_sram_buff_w12[116],loc_sram_buff_w12[117],loc_sram_buff_w12[118],loc_sram_buff_w12[119],loc_sram_buff_w12[120],loc_sram_buff_w12[121],loc_sram_buff_w12[122],loc_sram_buff_w12[123],loc_sram_buff_w12[124],loc_sram_buff_w12[125],loc_sram_buff_w12[126],loc_sram_buff_w12[127],loc_sram_buff_w12[128],loc_sram_buff_w12[129],loc_sram_buff_w12[130],loc_sram_buff_w12[131],loc_sram_buff_w12[132],loc_sram_buff_w12[133],loc_sram_buff_w12[134],loc_sram_buff_w12[135],loc_sram_buff_w12[136],loc_sram_buff_w12[137],loc_sram_buff_w12[138],loc_sram_buff_w12[139],loc_sram_buff_w12[140],loc_sram_buff_w12[141],loc_sram_buff_w12[142],loc_sram_buff_w12[143],loc_sram_buff_w12[144],loc_sram_buff_w12[145],loc_sram_buff_w12[146],loc_sram_buff_w12[147],loc_sram_buff_w12[148],loc_sram_buff_w12[149],loc_sram_buff_w12[150],loc_sram_buff_w12[151],loc_sram_buff_w12[152],loc_sram_buff_w12[153],loc_sram_buff_w12[154],loc_sram_buff_w12[155],loc_sram_buff_w12[156],loc_sram_buff_w12[157],loc_sram_buff_w12[158],loc_sram_buff_w12[159],loc_sram_buff_w12[160],loc_sram_buff_w12[161],loc_sram_buff_w12[162],loc_sram_buff_w12[163],loc_sram_buff_w12[164],loc_sram_buff_w12[165],loc_sram_buff_w12[166],loc_sram_buff_w12[167],loc_sram_buff_w12[168],loc_sram_buff_w12[169],loc_sram_buff_w12[170],loc_sram_buff_w12[171],loc_sram_buff_w12[172],loc_sram_buff_w12[173],loc_sram_buff_w12[174],loc_sram_buff_w12[175],loc_sram_buff_w12[176],loc_sram_buff_w12[177],loc_sram_buff_w12[178],loc_sram_buff_w12[179],loc_sram_buff_w12[180],loc_sram_buff_w12[181],loc_sram_buff_w12[182],loc_sram_buff_w12[183],loc_sram_buff_w12[184],loc_sram_buff_w12[185],loc_sram_buff_w12[186],loc_sram_buff_w12[187],loc_sram_buff_w12[188],loc_sram_buff_w12[189],loc_sram_buff_w12[190],loc_sram_buff_w12[191],loc_sram_buff_w12[192],loc_sram_buff_w12[193],loc_sram_buff_w12[194],loc_sram_buff_w12[195],loc_sram_buff_w12[196],loc_sram_buff_w12[197],loc_sram_buff_w12[198],loc_sram_buff_w12[199],loc_sram_buff_w12[200],loc_sram_buff_w12[201],loc_sram_buff_w12[202],loc_sram_buff_w12[203],loc_sram_buff_w12[204],loc_sram_buff_w12[205],loc_sram_buff_w12[206],loc_sram_buff_w12[207],loc_sram_buff_w12[208],loc_sram_buff_w12[209],loc_sram_buff_w12[210],loc_sram_buff_w12[211],loc_sram_buff_w12[212],loc_sram_buff_w12[213],loc_sram_buff_w12[214],loc_sram_buff_w12[215],loc_sram_buff_w12[216],loc_sram_buff_w12[217],loc_sram_buff_w12[218],loc_sram_buff_w12[219],loc_sram_buff_w12[220],loc_sram_buff_w12[221],loc_sram_buff_w12[222],loc_sram_buff_w12[223],loc_sram_buff_w12[224],loc_sram_buff_w12[225],loc_sram_buff_w12[226],loc_sram_buff_w12[227],loc_sram_buff_w12[228],loc_sram_buff_w12[229],loc_sram_buff_w12[230],loc_sram_buff_w12[231],loc_sram_buff_w12[232],loc_sram_buff_w12[233],loc_sram_buff_w12[234],loc_sram_buff_w12[235],loc_sram_buff_w12[236],loc_sram_buff_w12[237],loc_sram_buff_w12[238],loc_sram_buff_w12[239],loc_sram_buff_w12[240],loc_sram_buff_w12[241],loc_sram_buff_w12[242],loc_sram_buff_w12[243],loc_sram_buff_w12[244],loc_sram_buff_w12[245],loc_sram_buff_w12[246],loc_sram_buff_w12[247],loc_sram_buff_w12[248],loc_sram_buff_w12[249],loc_sram_buff_w12[250],loc_sram_buff_w12[251],loc_sram_buff_w12[252],loc_sram_buff_w12[253],loc_sram_buff_w12[254],loc_sram_buff_w12[255]} = loc_sram_rdata12;
	{loc_sram_buff_w13[0],loc_sram_buff_w13[1],loc_sram_buff_w13[2],loc_sram_buff_w13[3],loc_sram_buff_w13[4],loc_sram_buff_w13[5],loc_sram_buff_w13[6],loc_sram_buff_w13[7],loc_sram_buff_w13[8],loc_sram_buff_w13[9],loc_sram_buff_w13[10],loc_sram_buff_w13[11],loc_sram_buff_w13[12],loc_sram_buff_w13[13],loc_sram_buff_w13[14],loc_sram_buff_w13[15],loc_sram_buff_w13[16],loc_sram_buff_w13[17],loc_sram_buff_w13[18],loc_sram_buff_w13[19],loc_sram_buff_w13[20],loc_sram_buff_w13[21],loc_sram_buff_w13[22],loc_sram_buff_w13[23],loc_sram_buff_w13[24],loc_sram_buff_w13[25],loc_sram_buff_w13[26],loc_sram_buff_w13[27],loc_sram_buff_w13[28],loc_sram_buff_w13[29],loc_sram_buff_w13[30],loc_sram_buff_w13[31],loc_sram_buff_w13[32],loc_sram_buff_w13[33],loc_sram_buff_w13[34],loc_sram_buff_w13[35],loc_sram_buff_w13[36],loc_sram_buff_w13[37],loc_sram_buff_w13[38],loc_sram_buff_w13[39],loc_sram_buff_w13[40],loc_sram_buff_w13[41],loc_sram_buff_w13[42],loc_sram_buff_w13[43],loc_sram_buff_w13[44],loc_sram_buff_w13[45],loc_sram_buff_w13[46],loc_sram_buff_w13[47],loc_sram_buff_w13[48],loc_sram_buff_w13[49],loc_sram_buff_w13[50],loc_sram_buff_w13[51],loc_sram_buff_w13[52],loc_sram_buff_w13[53],loc_sram_buff_w13[54],loc_sram_buff_w13[55],loc_sram_buff_w13[56],loc_sram_buff_w13[57],loc_sram_buff_w13[58],loc_sram_buff_w13[59],loc_sram_buff_w13[60],loc_sram_buff_w13[61],loc_sram_buff_w13[62],loc_sram_buff_w13[63],loc_sram_buff_w13[64],loc_sram_buff_w13[65],loc_sram_buff_w13[66],loc_sram_buff_w13[67],loc_sram_buff_w13[68],loc_sram_buff_w13[69],loc_sram_buff_w13[70],loc_sram_buff_w13[71],loc_sram_buff_w13[72],loc_sram_buff_w13[73],loc_sram_buff_w13[74],loc_sram_buff_w13[75],loc_sram_buff_w13[76],loc_sram_buff_w13[77],loc_sram_buff_w13[78],loc_sram_buff_w13[79],loc_sram_buff_w13[80],loc_sram_buff_w13[81],loc_sram_buff_w13[82],loc_sram_buff_w13[83],loc_sram_buff_w13[84],loc_sram_buff_w13[85],loc_sram_buff_w13[86],loc_sram_buff_w13[87],loc_sram_buff_w13[88],loc_sram_buff_w13[89],loc_sram_buff_w13[90],loc_sram_buff_w13[91],loc_sram_buff_w13[92],loc_sram_buff_w13[93],loc_sram_buff_w13[94],loc_sram_buff_w13[95],loc_sram_buff_w13[96],loc_sram_buff_w13[97],loc_sram_buff_w13[98],loc_sram_buff_w13[99],loc_sram_buff_w13[100],loc_sram_buff_w13[101],loc_sram_buff_w13[102],loc_sram_buff_w13[103],loc_sram_buff_w13[104],loc_sram_buff_w13[105],loc_sram_buff_w13[106],loc_sram_buff_w13[107],loc_sram_buff_w13[108],loc_sram_buff_w13[109],loc_sram_buff_w13[110],loc_sram_buff_w13[111],loc_sram_buff_w13[112],loc_sram_buff_w13[113],loc_sram_buff_w13[114],loc_sram_buff_w13[115],loc_sram_buff_w13[116],loc_sram_buff_w13[117],loc_sram_buff_w13[118],loc_sram_buff_w13[119],loc_sram_buff_w13[120],loc_sram_buff_w13[121],loc_sram_buff_w13[122],loc_sram_buff_w13[123],loc_sram_buff_w13[124],loc_sram_buff_w13[125],loc_sram_buff_w13[126],loc_sram_buff_w13[127],loc_sram_buff_w13[128],loc_sram_buff_w13[129],loc_sram_buff_w13[130],loc_sram_buff_w13[131],loc_sram_buff_w13[132],loc_sram_buff_w13[133],loc_sram_buff_w13[134],loc_sram_buff_w13[135],loc_sram_buff_w13[136],loc_sram_buff_w13[137],loc_sram_buff_w13[138],loc_sram_buff_w13[139],loc_sram_buff_w13[140],loc_sram_buff_w13[141],loc_sram_buff_w13[142],loc_sram_buff_w13[143],loc_sram_buff_w13[144],loc_sram_buff_w13[145],loc_sram_buff_w13[146],loc_sram_buff_w13[147],loc_sram_buff_w13[148],loc_sram_buff_w13[149],loc_sram_buff_w13[150],loc_sram_buff_w13[151],loc_sram_buff_w13[152],loc_sram_buff_w13[153],loc_sram_buff_w13[154],loc_sram_buff_w13[155],loc_sram_buff_w13[156],loc_sram_buff_w13[157],loc_sram_buff_w13[158],loc_sram_buff_w13[159],loc_sram_buff_w13[160],loc_sram_buff_w13[161],loc_sram_buff_w13[162],loc_sram_buff_w13[163],loc_sram_buff_w13[164],loc_sram_buff_w13[165],loc_sram_buff_w13[166],loc_sram_buff_w13[167],loc_sram_buff_w13[168],loc_sram_buff_w13[169],loc_sram_buff_w13[170],loc_sram_buff_w13[171],loc_sram_buff_w13[172],loc_sram_buff_w13[173],loc_sram_buff_w13[174],loc_sram_buff_w13[175],loc_sram_buff_w13[176],loc_sram_buff_w13[177],loc_sram_buff_w13[178],loc_sram_buff_w13[179],loc_sram_buff_w13[180],loc_sram_buff_w13[181],loc_sram_buff_w13[182],loc_sram_buff_w13[183],loc_sram_buff_w13[184],loc_sram_buff_w13[185],loc_sram_buff_w13[186],loc_sram_buff_w13[187],loc_sram_buff_w13[188],loc_sram_buff_w13[189],loc_sram_buff_w13[190],loc_sram_buff_w13[191],loc_sram_buff_w13[192],loc_sram_buff_w13[193],loc_sram_buff_w13[194],loc_sram_buff_w13[195],loc_sram_buff_w13[196],loc_sram_buff_w13[197],loc_sram_buff_w13[198],loc_sram_buff_w13[199],loc_sram_buff_w13[200],loc_sram_buff_w13[201],loc_sram_buff_w13[202],loc_sram_buff_w13[203],loc_sram_buff_w13[204],loc_sram_buff_w13[205],loc_sram_buff_w13[206],loc_sram_buff_w13[207],loc_sram_buff_w13[208],loc_sram_buff_w13[209],loc_sram_buff_w13[210],loc_sram_buff_w13[211],loc_sram_buff_w13[212],loc_sram_buff_w13[213],loc_sram_buff_w13[214],loc_sram_buff_w13[215],loc_sram_buff_w13[216],loc_sram_buff_w13[217],loc_sram_buff_w13[218],loc_sram_buff_w13[219],loc_sram_buff_w13[220],loc_sram_buff_w13[221],loc_sram_buff_w13[222],loc_sram_buff_w13[223],loc_sram_buff_w13[224],loc_sram_buff_w13[225],loc_sram_buff_w13[226],loc_sram_buff_w13[227],loc_sram_buff_w13[228],loc_sram_buff_w13[229],loc_sram_buff_w13[230],loc_sram_buff_w13[231],loc_sram_buff_w13[232],loc_sram_buff_w13[233],loc_sram_buff_w13[234],loc_sram_buff_w13[235],loc_sram_buff_w13[236],loc_sram_buff_w13[237],loc_sram_buff_w13[238],loc_sram_buff_w13[239],loc_sram_buff_w13[240],loc_sram_buff_w13[241],loc_sram_buff_w13[242],loc_sram_buff_w13[243],loc_sram_buff_w13[244],loc_sram_buff_w13[245],loc_sram_buff_w13[246],loc_sram_buff_w13[247],loc_sram_buff_w13[248],loc_sram_buff_w13[249],loc_sram_buff_w13[250],loc_sram_buff_w13[251],loc_sram_buff_w13[252],loc_sram_buff_w13[253],loc_sram_buff_w13[254],loc_sram_buff_w13[255]} = loc_sram_rdata13;
	{loc_sram_buff_w14[0],loc_sram_buff_w14[1],loc_sram_buff_w14[2],loc_sram_buff_w14[3],loc_sram_buff_w14[4],loc_sram_buff_w14[5],loc_sram_buff_w14[6],loc_sram_buff_w14[7],loc_sram_buff_w14[8],loc_sram_buff_w14[9],loc_sram_buff_w14[10],loc_sram_buff_w14[11],loc_sram_buff_w14[12],loc_sram_buff_w14[13],loc_sram_buff_w14[14],loc_sram_buff_w14[15],loc_sram_buff_w14[16],loc_sram_buff_w14[17],loc_sram_buff_w14[18],loc_sram_buff_w14[19],loc_sram_buff_w14[20],loc_sram_buff_w14[21],loc_sram_buff_w14[22],loc_sram_buff_w14[23],loc_sram_buff_w14[24],loc_sram_buff_w14[25],loc_sram_buff_w14[26],loc_sram_buff_w14[27],loc_sram_buff_w14[28],loc_sram_buff_w14[29],loc_sram_buff_w14[30],loc_sram_buff_w14[31],loc_sram_buff_w14[32],loc_sram_buff_w14[33],loc_sram_buff_w14[34],loc_sram_buff_w14[35],loc_sram_buff_w14[36],loc_sram_buff_w14[37],loc_sram_buff_w14[38],loc_sram_buff_w14[39],loc_sram_buff_w14[40],loc_sram_buff_w14[41],loc_sram_buff_w14[42],loc_sram_buff_w14[43],loc_sram_buff_w14[44],loc_sram_buff_w14[45],loc_sram_buff_w14[46],loc_sram_buff_w14[47],loc_sram_buff_w14[48],loc_sram_buff_w14[49],loc_sram_buff_w14[50],loc_sram_buff_w14[51],loc_sram_buff_w14[52],loc_sram_buff_w14[53],loc_sram_buff_w14[54],loc_sram_buff_w14[55],loc_sram_buff_w14[56],loc_sram_buff_w14[57],loc_sram_buff_w14[58],loc_sram_buff_w14[59],loc_sram_buff_w14[60],loc_sram_buff_w14[61],loc_sram_buff_w14[62],loc_sram_buff_w14[63],loc_sram_buff_w14[64],loc_sram_buff_w14[65],loc_sram_buff_w14[66],loc_sram_buff_w14[67],loc_sram_buff_w14[68],loc_sram_buff_w14[69],loc_sram_buff_w14[70],loc_sram_buff_w14[71],loc_sram_buff_w14[72],loc_sram_buff_w14[73],loc_sram_buff_w14[74],loc_sram_buff_w14[75],loc_sram_buff_w14[76],loc_sram_buff_w14[77],loc_sram_buff_w14[78],loc_sram_buff_w14[79],loc_sram_buff_w14[80],loc_sram_buff_w14[81],loc_sram_buff_w14[82],loc_sram_buff_w14[83],loc_sram_buff_w14[84],loc_sram_buff_w14[85],loc_sram_buff_w14[86],loc_sram_buff_w14[87],loc_sram_buff_w14[88],loc_sram_buff_w14[89],loc_sram_buff_w14[90],loc_sram_buff_w14[91],loc_sram_buff_w14[92],loc_sram_buff_w14[93],loc_sram_buff_w14[94],loc_sram_buff_w14[95],loc_sram_buff_w14[96],loc_sram_buff_w14[97],loc_sram_buff_w14[98],loc_sram_buff_w14[99],loc_sram_buff_w14[100],loc_sram_buff_w14[101],loc_sram_buff_w14[102],loc_sram_buff_w14[103],loc_sram_buff_w14[104],loc_sram_buff_w14[105],loc_sram_buff_w14[106],loc_sram_buff_w14[107],loc_sram_buff_w14[108],loc_sram_buff_w14[109],loc_sram_buff_w14[110],loc_sram_buff_w14[111],loc_sram_buff_w14[112],loc_sram_buff_w14[113],loc_sram_buff_w14[114],loc_sram_buff_w14[115],loc_sram_buff_w14[116],loc_sram_buff_w14[117],loc_sram_buff_w14[118],loc_sram_buff_w14[119],loc_sram_buff_w14[120],loc_sram_buff_w14[121],loc_sram_buff_w14[122],loc_sram_buff_w14[123],loc_sram_buff_w14[124],loc_sram_buff_w14[125],loc_sram_buff_w14[126],loc_sram_buff_w14[127],loc_sram_buff_w14[128],loc_sram_buff_w14[129],loc_sram_buff_w14[130],loc_sram_buff_w14[131],loc_sram_buff_w14[132],loc_sram_buff_w14[133],loc_sram_buff_w14[134],loc_sram_buff_w14[135],loc_sram_buff_w14[136],loc_sram_buff_w14[137],loc_sram_buff_w14[138],loc_sram_buff_w14[139],loc_sram_buff_w14[140],loc_sram_buff_w14[141],loc_sram_buff_w14[142],loc_sram_buff_w14[143],loc_sram_buff_w14[144],loc_sram_buff_w14[145],loc_sram_buff_w14[146],loc_sram_buff_w14[147],loc_sram_buff_w14[148],loc_sram_buff_w14[149],loc_sram_buff_w14[150],loc_sram_buff_w14[151],loc_sram_buff_w14[152],loc_sram_buff_w14[153],loc_sram_buff_w14[154],loc_sram_buff_w14[155],loc_sram_buff_w14[156],loc_sram_buff_w14[157],loc_sram_buff_w14[158],loc_sram_buff_w14[159],loc_sram_buff_w14[160],loc_sram_buff_w14[161],loc_sram_buff_w14[162],loc_sram_buff_w14[163],loc_sram_buff_w14[164],loc_sram_buff_w14[165],loc_sram_buff_w14[166],loc_sram_buff_w14[167],loc_sram_buff_w14[168],loc_sram_buff_w14[169],loc_sram_buff_w14[170],loc_sram_buff_w14[171],loc_sram_buff_w14[172],loc_sram_buff_w14[173],loc_sram_buff_w14[174],loc_sram_buff_w14[175],loc_sram_buff_w14[176],loc_sram_buff_w14[177],loc_sram_buff_w14[178],loc_sram_buff_w14[179],loc_sram_buff_w14[180],loc_sram_buff_w14[181],loc_sram_buff_w14[182],loc_sram_buff_w14[183],loc_sram_buff_w14[184],loc_sram_buff_w14[185],loc_sram_buff_w14[186],loc_sram_buff_w14[187],loc_sram_buff_w14[188],loc_sram_buff_w14[189],loc_sram_buff_w14[190],loc_sram_buff_w14[191],loc_sram_buff_w14[192],loc_sram_buff_w14[193],loc_sram_buff_w14[194],loc_sram_buff_w14[195],loc_sram_buff_w14[196],loc_sram_buff_w14[197],loc_sram_buff_w14[198],loc_sram_buff_w14[199],loc_sram_buff_w14[200],loc_sram_buff_w14[201],loc_sram_buff_w14[202],loc_sram_buff_w14[203],loc_sram_buff_w14[204],loc_sram_buff_w14[205],loc_sram_buff_w14[206],loc_sram_buff_w14[207],loc_sram_buff_w14[208],loc_sram_buff_w14[209],loc_sram_buff_w14[210],loc_sram_buff_w14[211],loc_sram_buff_w14[212],loc_sram_buff_w14[213],loc_sram_buff_w14[214],loc_sram_buff_w14[215],loc_sram_buff_w14[216],loc_sram_buff_w14[217],loc_sram_buff_w14[218],loc_sram_buff_w14[219],loc_sram_buff_w14[220],loc_sram_buff_w14[221],loc_sram_buff_w14[222],loc_sram_buff_w14[223],loc_sram_buff_w14[224],loc_sram_buff_w14[225],loc_sram_buff_w14[226],loc_sram_buff_w14[227],loc_sram_buff_w14[228],loc_sram_buff_w14[229],loc_sram_buff_w14[230],loc_sram_buff_w14[231],loc_sram_buff_w14[232],loc_sram_buff_w14[233],loc_sram_buff_w14[234],loc_sram_buff_w14[235],loc_sram_buff_w14[236],loc_sram_buff_w14[237],loc_sram_buff_w14[238],loc_sram_buff_w14[239],loc_sram_buff_w14[240],loc_sram_buff_w14[241],loc_sram_buff_w14[242],loc_sram_buff_w14[243],loc_sram_buff_w14[244],loc_sram_buff_w14[245],loc_sram_buff_w14[246],loc_sram_buff_w14[247],loc_sram_buff_w14[248],loc_sram_buff_w14[249],loc_sram_buff_w14[250],loc_sram_buff_w14[251],loc_sram_buff_w14[252],loc_sram_buff_w14[253],loc_sram_buff_w14[254],loc_sram_buff_w14[255]} = loc_sram_rdata14;
	{loc_sram_buff_w15[0],loc_sram_buff_w15[1],loc_sram_buff_w15[2],loc_sram_buff_w15[3],loc_sram_buff_w15[4],loc_sram_buff_w15[5],loc_sram_buff_w15[6],loc_sram_buff_w15[7],loc_sram_buff_w15[8],loc_sram_buff_w15[9],loc_sram_buff_w15[10],loc_sram_buff_w15[11],loc_sram_buff_w15[12],loc_sram_buff_w15[13],loc_sram_buff_w15[14],loc_sram_buff_w15[15],loc_sram_buff_w15[16],loc_sram_buff_w15[17],loc_sram_buff_w15[18],loc_sram_buff_w15[19],loc_sram_buff_w15[20],loc_sram_buff_w15[21],loc_sram_buff_w15[22],loc_sram_buff_w15[23],loc_sram_buff_w15[24],loc_sram_buff_w15[25],loc_sram_buff_w15[26],loc_sram_buff_w15[27],loc_sram_buff_w15[28],loc_sram_buff_w15[29],loc_sram_buff_w15[30],loc_sram_buff_w15[31],loc_sram_buff_w15[32],loc_sram_buff_w15[33],loc_sram_buff_w15[34],loc_sram_buff_w15[35],loc_sram_buff_w15[36],loc_sram_buff_w15[37],loc_sram_buff_w15[38],loc_sram_buff_w15[39],loc_sram_buff_w15[40],loc_sram_buff_w15[41],loc_sram_buff_w15[42],loc_sram_buff_w15[43],loc_sram_buff_w15[44],loc_sram_buff_w15[45],loc_sram_buff_w15[46],loc_sram_buff_w15[47],loc_sram_buff_w15[48],loc_sram_buff_w15[49],loc_sram_buff_w15[50],loc_sram_buff_w15[51],loc_sram_buff_w15[52],loc_sram_buff_w15[53],loc_sram_buff_w15[54],loc_sram_buff_w15[55],loc_sram_buff_w15[56],loc_sram_buff_w15[57],loc_sram_buff_w15[58],loc_sram_buff_w15[59],loc_sram_buff_w15[60],loc_sram_buff_w15[61],loc_sram_buff_w15[62],loc_sram_buff_w15[63],loc_sram_buff_w15[64],loc_sram_buff_w15[65],loc_sram_buff_w15[66],loc_sram_buff_w15[67],loc_sram_buff_w15[68],loc_sram_buff_w15[69],loc_sram_buff_w15[70],loc_sram_buff_w15[71],loc_sram_buff_w15[72],loc_sram_buff_w15[73],loc_sram_buff_w15[74],loc_sram_buff_w15[75],loc_sram_buff_w15[76],loc_sram_buff_w15[77],loc_sram_buff_w15[78],loc_sram_buff_w15[79],loc_sram_buff_w15[80],loc_sram_buff_w15[81],loc_sram_buff_w15[82],loc_sram_buff_w15[83],loc_sram_buff_w15[84],loc_sram_buff_w15[85],loc_sram_buff_w15[86],loc_sram_buff_w15[87],loc_sram_buff_w15[88],loc_sram_buff_w15[89],loc_sram_buff_w15[90],loc_sram_buff_w15[91],loc_sram_buff_w15[92],loc_sram_buff_w15[93],loc_sram_buff_w15[94],loc_sram_buff_w15[95],loc_sram_buff_w15[96],loc_sram_buff_w15[97],loc_sram_buff_w15[98],loc_sram_buff_w15[99],loc_sram_buff_w15[100],loc_sram_buff_w15[101],loc_sram_buff_w15[102],loc_sram_buff_w15[103],loc_sram_buff_w15[104],loc_sram_buff_w15[105],loc_sram_buff_w15[106],loc_sram_buff_w15[107],loc_sram_buff_w15[108],loc_sram_buff_w15[109],loc_sram_buff_w15[110],loc_sram_buff_w15[111],loc_sram_buff_w15[112],loc_sram_buff_w15[113],loc_sram_buff_w15[114],loc_sram_buff_w15[115],loc_sram_buff_w15[116],loc_sram_buff_w15[117],loc_sram_buff_w15[118],loc_sram_buff_w15[119],loc_sram_buff_w15[120],loc_sram_buff_w15[121],loc_sram_buff_w15[122],loc_sram_buff_w15[123],loc_sram_buff_w15[124],loc_sram_buff_w15[125],loc_sram_buff_w15[126],loc_sram_buff_w15[127],loc_sram_buff_w15[128],loc_sram_buff_w15[129],loc_sram_buff_w15[130],loc_sram_buff_w15[131],loc_sram_buff_w15[132],loc_sram_buff_w15[133],loc_sram_buff_w15[134],loc_sram_buff_w15[135],loc_sram_buff_w15[136],loc_sram_buff_w15[137],loc_sram_buff_w15[138],loc_sram_buff_w15[139],loc_sram_buff_w15[140],loc_sram_buff_w15[141],loc_sram_buff_w15[142],loc_sram_buff_w15[143],loc_sram_buff_w15[144],loc_sram_buff_w15[145],loc_sram_buff_w15[146],loc_sram_buff_w15[147],loc_sram_buff_w15[148],loc_sram_buff_w15[149],loc_sram_buff_w15[150],loc_sram_buff_w15[151],loc_sram_buff_w15[152],loc_sram_buff_w15[153],loc_sram_buff_w15[154],loc_sram_buff_w15[155],loc_sram_buff_w15[156],loc_sram_buff_w15[157],loc_sram_buff_w15[158],loc_sram_buff_w15[159],loc_sram_buff_w15[160],loc_sram_buff_w15[161],loc_sram_buff_w15[162],loc_sram_buff_w15[163],loc_sram_buff_w15[164],loc_sram_buff_w15[165],loc_sram_buff_w15[166],loc_sram_buff_w15[167],loc_sram_buff_w15[168],loc_sram_buff_w15[169],loc_sram_buff_w15[170],loc_sram_buff_w15[171],loc_sram_buff_w15[172],loc_sram_buff_w15[173],loc_sram_buff_w15[174],loc_sram_buff_w15[175],loc_sram_buff_w15[176],loc_sram_buff_w15[177],loc_sram_buff_w15[178],loc_sram_buff_w15[179],loc_sram_buff_w15[180],loc_sram_buff_w15[181],loc_sram_buff_w15[182],loc_sram_buff_w15[183],loc_sram_buff_w15[184],loc_sram_buff_w15[185],loc_sram_buff_w15[186],loc_sram_buff_w15[187],loc_sram_buff_w15[188],loc_sram_buff_w15[189],loc_sram_buff_w15[190],loc_sram_buff_w15[191],loc_sram_buff_w15[192],loc_sram_buff_w15[193],loc_sram_buff_w15[194],loc_sram_buff_w15[195],loc_sram_buff_w15[196],loc_sram_buff_w15[197],loc_sram_buff_w15[198],loc_sram_buff_w15[199],loc_sram_buff_w15[200],loc_sram_buff_w15[201],loc_sram_buff_w15[202],loc_sram_buff_w15[203],loc_sram_buff_w15[204],loc_sram_buff_w15[205],loc_sram_buff_w15[206],loc_sram_buff_w15[207],loc_sram_buff_w15[208],loc_sram_buff_w15[209],loc_sram_buff_w15[210],loc_sram_buff_w15[211],loc_sram_buff_w15[212],loc_sram_buff_w15[213],loc_sram_buff_w15[214],loc_sram_buff_w15[215],loc_sram_buff_w15[216],loc_sram_buff_w15[217],loc_sram_buff_w15[218],loc_sram_buff_w15[219],loc_sram_buff_w15[220],loc_sram_buff_w15[221],loc_sram_buff_w15[222],loc_sram_buff_w15[223],loc_sram_buff_w15[224],loc_sram_buff_w15[225],loc_sram_buff_w15[226],loc_sram_buff_w15[227],loc_sram_buff_w15[228],loc_sram_buff_w15[229],loc_sram_buff_w15[230],loc_sram_buff_w15[231],loc_sram_buff_w15[232],loc_sram_buff_w15[233],loc_sram_buff_w15[234],loc_sram_buff_w15[235],loc_sram_buff_w15[236],loc_sram_buff_w15[237],loc_sram_buff_w15[238],loc_sram_buff_w15[239],loc_sram_buff_w15[240],loc_sram_buff_w15[241],loc_sram_buff_w15[242],loc_sram_buff_w15[243],loc_sram_buff_w15[244],loc_sram_buff_w15[245],loc_sram_buff_w15[246],loc_sram_buff_w15[247],loc_sram_buff_w15[248],loc_sram_buff_w15[249],loc_sram_buff_w15[250],loc_sram_buff_w15[251],loc_sram_buff_w15[252],loc_sram_buff_w15[253],loc_sram_buff_w15[254],loc_sram_buff_w15[255]} = loc_sram_rdata15;

		
	loc_rdata_buff[1023:1020] = ({4{loc_sram_buff_w0[0][4]}} & loc_sram_buff_w0[0][3:0]) | ({4{loc_sram_buff_w1[0][4]}} & loc_sram_buff_w1[0][3:0]) | ({4{loc_sram_buff_w2[0][4]}} & loc_sram_buff_w2[0][3:0]) | ({4{loc_sram_buff_w3[0][4]}} & loc_sram_buff_w3[0][3:0]) | ({4{loc_sram_buff_w4[0][4]}} & loc_sram_buff_w4[0][3:0]) | ({4{loc_sram_buff_w5[0][4]}} & loc_sram_buff_w5[0][3:0]) | ({4{loc_sram_buff_w6[0][4]}} & loc_sram_buff_w6[0][3:0]) | ({4{loc_sram_buff_w7[0][4]}} & loc_sram_buff_w7[0][3:0]) | ({4{loc_sram_buff_w8[0][4]}} & loc_sram_buff_w8[0][3:0]) | ({4{loc_sram_buff_w9[0][4]}} & loc_sram_buff_w9[0][3:0]) | ({4{loc_sram_buff_w10[0][4]}} & loc_sram_buff_w10[0][3:0]) | ({4{loc_sram_buff_w11[0][4]}} & loc_sram_buff_w11[0][3:0]) | ({4{loc_sram_buff_w12[0][4]}} & loc_sram_buff_w12[0][3:0]) | ({4{loc_sram_buff_w13[0][4]}} & loc_sram_buff_w13[0][3:0]) | ({4{loc_sram_buff_w14[0][4]}} & loc_sram_buff_w14[0][3:0]) | ({4{loc_sram_buff_w15[0][4]}} & loc_sram_buff_w15[0][3:0]);
	loc_rdata_buff[1019:1016] = ({4{loc_sram_buff_w0[1][4]}} & loc_sram_buff_w0[1][3:0]) | ({4{loc_sram_buff_w1[1][4]}} & loc_sram_buff_w1[1][3:0]) | ({4{loc_sram_buff_w2[1][4]}} & loc_sram_buff_w2[1][3:0]) | ({4{loc_sram_buff_w3[1][4]}} & loc_sram_buff_w3[1][3:0]) | ({4{loc_sram_buff_w4[1][4]}} & loc_sram_buff_w4[1][3:0]) | ({4{loc_sram_buff_w5[1][4]}} & loc_sram_buff_w5[1][3:0]) | ({4{loc_sram_buff_w6[1][4]}} & loc_sram_buff_w6[1][3:0]) | ({4{loc_sram_buff_w7[1][4]}} & loc_sram_buff_w7[1][3:0]) | ({4{loc_sram_buff_w8[1][4]}} & loc_sram_buff_w8[1][3:0]) | ({4{loc_sram_buff_w9[1][4]}} & loc_sram_buff_w9[1][3:0]) | ({4{loc_sram_buff_w10[1][4]}} & loc_sram_buff_w10[1][3:0]) | ({4{loc_sram_buff_w11[1][4]}} & loc_sram_buff_w11[1][3:0]) | ({4{loc_sram_buff_w12[1][4]}} & loc_sram_buff_w12[1][3:0]) | ({4{loc_sram_buff_w13[1][4]}} & loc_sram_buff_w13[1][3:0]) | ({4{loc_sram_buff_w14[1][4]}} & loc_sram_buff_w14[1][3:0]) | ({4{loc_sram_buff_w15[1][4]}} & loc_sram_buff_w15[1][3:0]);
	loc_rdata_buff[1015:1012] = ({4{loc_sram_buff_w0[2][4]}} & loc_sram_buff_w0[2][3:0]) | ({4{loc_sram_buff_w1[2][4]}} & loc_sram_buff_w1[2][3:0]) | ({4{loc_sram_buff_w2[2][4]}} & loc_sram_buff_w2[2][3:0]) | ({4{loc_sram_buff_w3[2][4]}} & loc_sram_buff_w3[2][3:0]) | ({4{loc_sram_buff_w4[2][4]}} & loc_sram_buff_w4[2][3:0]) | ({4{loc_sram_buff_w5[2][4]}} & loc_sram_buff_w5[2][3:0]) | ({4{loc_sram_buff_w6[2][4]}} & loc_sram_buff_w6[2][3:0]) | ({4{loc_sram_buff_w7[2][4]}} & loc_sram_buff_w7[2][3:0]) | ({4{loc_sram_buff_w8[2][4]}} & loc_sram_buff_w8[2][3:0]) | ({4{loc_sram_buff_w9[2][4]}} & loc_sram_buff_w9[2][3:0]) | ({4{loc_sram_buff_w10[2][4]}} & loc_sram_buff_w10[2][3:0]) | ({4{loc_sram_buff_w11[2][4]}} & loc_sram_buff_w11[2][3:0]) | ({4{loc_sram_buff_w12[2][4]}} & loc_sram_buff_w12[2][3:0]) | ({4{loc_sram_buff_w13[2][4]}} & loc_sram_buff_w13[2][3:0]) | ({4{loc_sram_buff_w14[2][4]}} & loc_sram_buff_w14[2][3:0]) | ({4{loc_sram_buff_w15[2][4]}} & loc_sram_buff_w15[2][3:0]);
	loc_rdata_buff[1011:1008] = ({4{loc_sram_buff_w0[3][4]}} & loc_sram_buff_w0[3][3:0]) | ({4{loc_sram_buff_w1[3][4]}} & loc_sram_buff_w1[3][3:0]) | ({4{loc_sram_buff_w2[3][4]}} & loc_sram_buff_w2[3][3:0]) | ({4{loc_sram_buff_w3[3][4]}} & loc_sram_buff_w3[3][3:0]) | ({4{loc_sram_buff_w4[3][4]}} & loc_sram_buff_w4[3][3:0]) | ({4{loc_sram_buff_w5[3][4]}} & loc_sram_buff_w5[3][3:0]) | ({4{loc_sram_buff_w6[3][4]}} & loc_sram_buff_w6[3][3:0]) | ({4{loc_sram_buff_w7[3][4]}} & loc_sram_buff_w7[3][3:0]) | ({4{loc_sram_buff_w8[3][4]}} & loc_sram_buff_w8[3][3:0]) | ({4{loc_sram_buff_w9[3][4]}} & loc_sram_buff_w9[3][3:0]) | ({4{loc_sram_buff_w10[3][4]}} & loc_sram_buff_w10[3][3:0]) | ({4{loc_sram_buff_w11[3][4]}} & loc_sram_buff_w11[3][3:0]) | ({4{loc_sram_buff_w12[3][4]}} & loc_sram_buff_w12[3][3:0]) | ({4{loc_sram_buff_w13[3][4]}} & loc_sram_buff_w13[3][3:0]) | ({4{loc_sram_buff_w14[3][4]}} & loc_sram_buff_w14[3][3:0]) | ({4{loc_sram_buff_w15[3][4]}} & loc_sram_buff_w15[3][3:0]);
	loc_rdata_buff[1007:1004] = ({4{loc_sram_buff_w0[4][4]}} & loc_sram_buff_w0[4][3:0]) | ({4{loc_sram_buff_w1[4][4]}} & loc_sram_buff_w1[4][3:0]) | ({4{loc_sram_buff_w2[4][4]}} & loc_sram_buff_w2[4][3:0]) | ({4{loc_sram_buff_w3[4][4]}} & loc_sram_buff_w3[4][3:0]) | ({4{loc_sram_buff_w4[4][4]}} & loc_sram_buff_w4[4][3:0]) | ({4{loc_sram_buff_w5[4][4]}} & loc_sram_buff_w5[4][3:0]) | ({4{loc_sram_buff_w6[4][4]}} & loc_sram_buff_w6[4][3:0]) | ({4{loc_sram_buff_w7[4][4]}} & loc_sram_buff_w7[4][3:0]) | ({4{loc_sram_buff_w8[4][4]}} & loc_sram_buff_w8[4][3:0]) | ({4{loc_sram_buff_w9[4][4]}} & loc_sram_buff_w9[4][3:0]) | ({4{loc_sram_buff_w10[4][4]}} & loc_sram_buff_w10[4][3:0]) | ({4{loc_sram_buff_w11[4][4]}} & loc_sram_buff_w11[4][3:0]) | ({4{loc_sram_buff_w12[4][4]}} & loc_sram_buff_w12[4][3:0]) | ({4{loc_sram_buff_w13[4][4]}} & loc_sram_buff_w13[4][3:0]) | ({4{loc_sram_buff_w14[4][4]}} & loc_sram_buff_w14[4][3:0]) | ({4{loc_sram_buff_w15[4][4]}} & loc_sram_buff_w15[4][3:0]);
	loc_rdata_buff[1003:1000] = ({4{loc_sram_buff_w0[5][4]}} & loc_sram_buff_w0[5][3:0]) | ({4{loc_sram_buff_w1[5][4]}} & loc_sram_buff_w1[5][3:0]) | ({4{loc_sram_buff_w2[5][4]}} & loc_sram_buff_w2[5][3:0]) | ({4{loc_sram_buff_w3[5][4]}} & loc_sram_buff_w3[5][3:0]) | ({4{loc_sram_buff_w4[5][4]}} & loc_sram_buff_w4[5][3:0]) | ({4{loc_sram_buff_w5[5][4]}} & loc_sram_buff_w5[5][3:0]) | ({4{loc_sram_buff_w6[5][4]}} & loc_sram_buff_w6[5][3:0]) | ({4{loc_sram_buff_w7[5][4]}} & loc_sram_buff_w7[5][3:0]) | ({4{loc_sram_buff_w8[5][4]}} & loc_sram_buff_w8[5][3:0]) | ({4{loc_sram_buff_w9[5][4]}} & loc_sram_buff_w9[5][3:0]) | ({4{loc_sram_buff_w10[5][4]}} & loc_sram_buff_w10[5][3:0]) | ({4{loc_sram_buff_w11[5][4]}} & loc_sram_buff_w11[5][3:0]) | ({4{loc_sram_buff_w12[5][4]}} & loc_sram_buff_w12[5][3:0]) | ({4{loc_sram_buff_w13[5][4]}} & loc_sram_buff_w13[5][3:0]) | ({4{loc_sram_buff_w14[5][4]}} & loc_sram_buff_w14[5][3:0]) | ({4{loc_sram_buff_w15[5][4]}} & loc_sram_buff_w15[5][3:0]);
	loc_rdata_buff[ 999: 996] = ({4{loc_sram_buff_w0[6][4]}} & loc_sram_buff_w0[6][3:0]) | ({4{loc_sram_buff_w1[6][4]}} & loc_sram_buff_w1[6][3:0]) | ({4{loc_sram_buff_w2[6][4]}} & loc_sram_buff_w2[6][3:0]) | ({4{loc_sram_buff_w3[6][4]}} & loc_sram_buff_w3[6][3:0]) | ({4{loc_sram_buff_w4[6][4]}} & loc_sram_buff_w4[6][3:0]) | ({4{loc_sram_buff_w5[6][4]}} & loc_sram_buff_w5[6][3:0]) | ({4{loc_sram_buff_w6[6][4]}} & loc_sram_buff_w6[6][3:0]) | ({4{loc_sram_buff_w7[6][4]}} & loc_sram_buff_w7[6][3:0]) | ({4{loc_sram_buff_w8[6][4]}} & loc_sram_buff_w8[6][3:0]) | ({4{loc_sram_buff_w9[6][4]}} & loc_sram_buff_w9[6][3:0]) | ({4{loc_sram_buff_w10[6][4]}} & loc_sram_buff_w10[6][3:0]) | ({4{loc_sram_buff_w11[6][4]}} & loc_sram_buff_w11[6][3:0]) | ({4{loc_sram_buff_w12[6][4]}} & loc_sram_buff_w12[6][3:0]) | ({4{loc_sram_buff_w13[6][4]}} & loc_sram_buff_w13[6][3:0]) | ({4{loc_sram_buff_w14[6][4]}} & loc_sram_buff_w14[6][3:0]) | ({4{loc_sram_buff_w15[6][4]}} & loc_sram_buff_w15[6][3:0]);
	loc_rdata_buff[ 995: 992] = ({4{loc_sram_buff_w0[7][4]}} & loc_sram_buff_w0[7][3:0]) | ({4{loc_sram_buff_w1[7][4]}} & loc_sram_buff_w1[7][3:0]) | ({4{loc_sram_buff_w2[7][4]}} & loc_sram_buff_w2[7][3:0]) | ({4{loc_sram_buff_w3[7][4]}} & loc_sram_buff_w3[7][3:0]) | ({4{loc_sram_buff_w4[7][4]}} & loc_sram_buff_w4[7][3:0]) | ({4{loc_sram_buff_w5[7][4]}} & loc_sram_buff_w5[7][3:0]) | ({4{loc_sram_buff_w6[7][4]}} & loc_sram_buff_w6[7][3:0]) | ({4{loc_sram_buff_w7[7][4]}} & loc_sram_buff_w7[7][3:0]) | ({4{loc_sram_buff_w8[7][4]}} & loc_sram_buff_w8[7][3:0]) | ({4{loc_sram_buff_w9[7][4]}} & loc_sram_buff_w9[7][3:0]) | ({4{loc_sram_buff_w10[7][4]}} & loc_sram_buff_w10[7][3:0]) | ({4{loc_sram_buff_w11[7][4]}} & loc_sram_buff_w11[7][3:0]) | ({4{loc_sram_buff_w12[7][4]}} & loc_sram_buff_w12[7][3:0]) | ({4{loc_sram_buff_w13[7][4]}} & loc_sram_buff_w13[7][3:0]) | ({4{loc_sram_buff_w14[7][4]}} & loc_sram_buff_w14[7][3:0]) | ({4{loc_sram_buff_w15[7][4]}} & loc_sram_buff_w15[7][3:0]);
	loc_rdata_buff[ 991: 988] = ({4{loc_sram_buff_w0[8][4]}} & loc_sram_buff_w0[8][3:0]) | ({4{loc_sram_buff_w1[8][4]}} & loc_sram_buff_w1[8][3:0]) | ({4{loc_sram_buff_w2[8][4]}} & loc_sram_buff_w2[8][3:0]) | ({4{loc_sram_buff_w3[8][4]}} & loc_sram_buff_w3[8][3:0]) | ({4{loc_sram_buff_w4[8][4]}} & loc_sram_buff_w4[8][3:0]) | ({4{loc_sram_buff_w5[8][4]}} & loc_sram_buff_w5[8][3:0]) | ({4{loc_sram_buff_w6[8][4]}} & loc_sram_buff_w6[8][3:0]) | ({4{loc_sram_buff_w7[8][4]}} & loc_sram_buff_w7[8][3:0]) | ({4{loc_sram_buff_w8[8][4]}} & loc_sram_buff_w8[8][3:0]) | ({4{loc_sram_buff_w9[8][4]}} & loc_sram_buff_w9[8][3:0]) | ({4{loc_sram_buff_w10[8][4]}} & loc_sram_buff_w10[8][3:0]) | ({4{loc_sram_buff_w11[8][4]}} & loc_sram_buff_w11[8][3:0]) | ({4{loc_sram_buff_w12[8][4]}} & loc_sram_buff_w12[8][3:0]) | ({4{loc_sram_buff_w13[8][4]}} & loc_sram_buff_w13[8][3:0]) | ({4{loc_sram_buff_w14[8][4]}} & loc_sram_buff_w14[8][3:0]) | ({4{loc_sram_buff_w15[8][4]}} & loc_sram_buff_w15[8][3:0]);
	loc_rdata_buff[ 987: 984] = ({4{loc_sram_buff_w0[9][4]}} & loc_sram_buff_w0[9][3:0]) | ({4{loc_sram_buff_w1[9][4]}} & loc_sram_buff_w1[9][3:0]) | ({4{loc_sram_buff_w2[9][4]}} & loc_sram_buff_w2[9][3:0]) | ({4{loc_sram_buff_w3[9][4]}} & loc_sram_buff_w3[9][3:0]) | ({4{loc_sram_buff_w4[9][4]}} & loc_sram_buff_w4[9][3:0]) | ({4{loc_sram_buff_w5[9][4]}} & loc_sram_buff_w5[9][3:0]) | ({4{loc_sram_buff_w6[9][4]}} & loc_sram_buff_w6[9][3:0]) | ({4{loc_sram_buff_w7[9][4]}} & loc_sram_buff_w7[9][3:0]) | ({4{loc_sram_buff_w8[9][4]}} & loc_sram_buff_w8[9][3:0]) | ({4{loc_sram_buff_w9[9][4]}} & loc_sram_buff_w9[9][3:0]) | ({4{loc_sram_buff_w10[9][4]}} & loc_sram_buff_w10[9][3:0]) | ({4{loc_sram_buff_w11[9][4]}} & loc_sram_buff_w11[9][3:0]) | ({4{loc_sram_buff_w12[9][4]}} & loc_sram_buff_w12[9][3:0]) | ({4{loc_sram_buff_w13[9][4]}} & loc_sram_buff_w13[9][3:0]) | ({4{loc_sram_buff_w14[9][4]}} & loc_sram_buff_w14[9][3:0]) | ({4{loc_sram_buff_w15[9][4]}} & loc_sram_buff_w15[9][3:0]);
	loc_rdata_buff[ 983: 980] = ({4{loc_sram_buff_w0[10][4]}} & loc_sram_buff_w0[10][3:0]) | ({4{loc_sram_buff_w1[10][4]}} & loc_sram_buff_w1[10][3:0]) | ({4{loc_sram_buff_w2[10][4]}} & loc_sram_buff_w2[10][3:0]) | ({4{loc_sram_buff_w3[10][4]}} & loc_sram_buff_w3[10][3:0]) | ({4{loc_sram_buff_w4[10][4]}} & loc_sram_buff_w4[10][3:0]) | ({4{loc_sram_buff_w5[10][4]}} & loc_sram_buff_w5[10][3:0]) | ({4{loc_sram_buff_w6[10][4]}} & loc_sram_buff_w6[10][3:0]) | ({4{loc_sram_buff_w7[10][4]}} & loc_sram_buff_w7[10][3:0]) | ({4{loc_sram_buff_w8[10][4]}} & loc_sram_buff_w8[10][3:0]) | ({4{loc_sram_buff_w9[10][4]}} & loc_sram_buff_w9[10][3:0]) | ({4{loc_sram_buff_w10[10][4]}} & loc_sram_buff_w10[10][3:0]) | ({4{loc_sram_buff_w11[10][4]}} & loc_sram_buff_w11[10][3:0]) | ({4{loc_sram_buff_w12[10][4]}} & loc_sram_buff_w12[10][3:0]) | ({4{loc_sram_buff_w13[10][4]}} & loc_sram_buff_w13[10][3:0]) | ({4{loc_sram_buff_w14[10][4]}} & loc_sram_buff_w14[10][3:0]) | ({4{loc_sram_buff_w15[10][4]}} & loc_sram_buff_w15[10][3:0]);
	loc_rdata_buff[ 979: 976] = ({4{loc_sram_buff_w0[11][4]}} & loc_sram_buff_w0[11][3:0]) | ({4{loc_sram_buff_w1[11][4]}} & loc_sram_buff_w1[11][3:0]) | ({4{loc_sram_buff_w2[11][4]}} & loc_sram_buff_w2[11][3:0]) | ({4{loc_sram_buff_w3[11][4]}} & loc_sram_buff_w3[11][3:0]) | ({4{loc_sram_buff_w4[11][4]}} & loc_sram_buff_w4[11][3:0]) | ({4{loc_sram_buff_w5[11][4]}} & loc_sram_buff_w5[11][3:0]) | ({4{loc_sram_buff_w6[11][4]}} & loc_sram_buff_w6[11][3:0]) | ({4{loc_sram_buff_w7[11][4]}} & loc_sram_buff_w7[11][3:0]) | ({4{loc_sram_buff_w8[11][4]}} & loc_sram_buff_w8[11][3:0]) | ({4{loc_sram_buff_w9[11][4]}} & loc_sram_buff_w9[11][3:0]) | ({4{loc_sram_buff_w10[11][4]}} & loc_sram_buff_w10[11][3:0]) | ({4{loc_sram_buff_w11[11][4]}} & loc_sram_buff_w11[11][3:0]) | ({4{loc_sram_buff_w12[11][4]}} & loc_sram_buff_w12[11][3:0]) | ({4{loc_sram_buff_w13[11][4]}} & loc_sram_buff_w13[11][3:0]) | ({4{loc_sram_buff_w14[11][4]}} & loc_sram_buff_w14[11][3:0]) | ({4{loc_sram_buff_w15[11][4]}} & loc_sram_buff_w15[11][3:0]);
	loc_rdata_buff[ 975: 972] = ({4{loc_sram_buff_w0[12][4]}} & loc_sram_buff_w0[12][3:0]) | ({4{loc_sram_buff_w1[12][4]}} & loc_sram_buff_w1[12][3:0]) | ({4{loc_sram_buff_w2[12][4]}} & loc_sram_buff_w2[12][3:0]) | ({4{loc_sram_buff_w3[12][4]}} & loc_sram_buff_w3[12][3:0]) | ({4{loc_sram_buff_w4[12][4]}} & loc_sram_buff_w4[12][3:0]) | ({4{loc_sram_buff_w5[12][4]}} & loc_sram_buff_w5[12][3:0]) | ({4{loc_sram_buff_w6[12][4]}} & loc_sram_buff_w6[12][3:0]) | ({4{loc_sram_buff_w7[12][4]}} & loc_sram_buff_w7[12][3:0]) | ({4{loc_sram_buff_w8[12][4]}} & loc_sram_buff_w8[12][3:0]) | ({4{loc_sram_buff_w9[12][4]}} & loc_sram_buff_w9[12][3:0]) | ({4{loc_sram_buff_w10[12][4]}} & loc_sram_buff_w10[12][3:0]) | ({4{loc_sram_buff_w11[12][4]}} & loc_sram_buff_w11[12][3:0]) | ({4{loc_sram_buff_w12[12][4]}} & loc_sram_buff_w12[12][3:0]) | ({4{loc_sram_buff_w13[12][4]}} & loc_sram_buff_w13[12][3:0]) | ({4{loc_sram_buff_w14[12][4]}} & loc_sram_buff_w14[12][3:0]) | ({4{loc_sram_buff_w15[12][4]}} & loc_sram_buff_w15[12][3:0]);
	loc_rdata_buff[ 971: 968] = ({4{loc_sram_buff_w0[13][4]}} & loc_sram_buff_w0[13][3:0]) | ({4{loc_sram_buff_w1[13][4]}} & loc_sram_buff_w1[13][3:0]) | ({4{loc_sram_buff_w2[13][4]}} & loc_sram_buff_w2[13][3:0]) | ({4{loc_sram_buff_w3[13][4]}} & loc_sram_buff_w3[13][3:0]) | ({4{loc_sram_buff_w4[13][4]}} & loc_sram_buff_w4[13][3:0]) | ({4{loc_sram_buff_w5[13][4]}} & loc_sram_buff_w5[13][3:0]) | ({4{loc_sram_buff_w6[13][4]}} & loc_sram_buff_w6[13][3:0]) | ({4{loc_sram_buff_w7[13][4]}} & loc_sram_buff_w7[13][3:0]) | ({4{loc_sram_buff_w8[13][4]}} & loc_sram_buff_w8[13][3:0]) | ({4{loc_sram_buff_w9[13][4]}} & loc_sram_buff_w9[13][3:0]) | ({4{loc_sram_buff_w10[13][4]}} & loc_sram_buff_w10[13][3:0]) | ({4{loc_sram_buff_w11[13][4]}} & loc_sram_buff_w11[13][3:0]) | ({4{loc_sram_buff_w12[13][4]}} & loc_sram_buff_w12[13][3:0]) | ({4{loc_sram_buff_w13[13][4]}} & loc_sram_buff_w13[13][3:0]) | ({4{loc_sram_buff_w14[13][4]}} & loc_sram_buff_w14[13][3:0]) | ({4{loc_sram_buff_w15[13][4]}} & loc_sram_buff_w15[13][3:0]);
	loc_rdata_buff[ 967: 964] = ({4{loc_sram_buff_w0[14][4]}} & loc_sram_buff_w0[14][3:0]) | ({4{loc_sram_buff_w1[14][4]}} & loc_sram_buff_w1[14][3:0]) | ({4{loc_sram_buff_w2[14][4]}} & loc_sram_buff_w2[14][3:0]) | ({4{loc_sram_buff_w3[14][4]}} & loc_sram_buff_w3[14][3:0]) | ({4{loc_sram_buff_w4[14][4]}} & loc_sram_buff_w4[14][3:0]) | ({4{loc_sram_buff_w5[14][4]}} & loc_sram_buff_w5[14][3:0]) | ({4{loc_sram_buff_w6[14][4]}} & loc_sram_buff_w6[14][3:0]) | ({4{loc_sram_buff_w7[14][4]}} & loc_sram_buff_w7[14][3:0]) | ({4{loc_sram_buff_w8[14][4]}} & loc_sram_buff_w8[14][3:0]) | ({4{loc_sram_buff_w9[14][4]}} & loc_sram_buff_w9[14][3:0]) | ({4{loc_sram_buff_w10[14][4]}} & loc_sram_buff_w10[14][3:0]) | ({4{loc_sram_buff_w11[14][4]}} & loc_sram_buff_w11[14][3:0]) | ({4{loc_sram_buff_w12[14][4]}} & loc_sram_buff_w12[14][3:0]) | ({4{loc_sram_buff_w13[14][4]}} & loc_sram_buff_w13[14][3:0]) | ({4{loc_sram_buff_w14[14][4]}} & loc_sram_buff_w14[14][3:0]) | ({4{loc_sram_buff_w15[14][4]}} & loc_sram_buff_w15[14][3:0]);
	loc_rdata_buff[ 963: 960] = ({4{loc_sram_buff_w0[15][4]}} & loc_sram_buff_w0[15][3:0]) | ({4{loc_sram_buff_w1[15][4]}} & loc_sram_buff_w1[15][3:0]) | ({4{loc_sram_buff_w2[15][4]}} & loc_sram_buff_w2[15][3:0]) | ({4{loc_sram_buff_w3[15][4]}} & loc_sram_buff_w3[15][3:0]) | ({4{loc_sram_buff_w4[15][4]}} & loc_sram_buff_w4[15][3:0]) | ({4{loc_sram_buff_w5[15][4]}} & loc_sram_buff_w5[15][3:0]) | ({4{loc_sram_buff_w6[15][4]}} & loc_sram_buff_w6[15][3:0]) | ({4{loc_sram_buff_w7[15][4]}} & loc_sram_buff_w7[15][3:0]) | ({4{loc_sram_buff_w8[15][4]}} & loc_sram_buff_w8[15][3:0]) | ({4{loc_sram_buff_w9[15][4]}} & loc_sram_buff_w9[15][3:0]) | ({4{loc_sram_buff_w10[15][4]}} & loc_sram_buff_w10[15][3:0]) | ({4{loc_sram_buff_w11[15][4]}} & loc_sram_buff_w11[15][3:0]) | ({4{loc_sram_buff_w12[15][4]}} & loc_sram_buff_w12[15][3:0]) | ({4{loc_sram_buff_w13[15][4]}} & loc_sram_buff_w13[15][3:0]) | ({4{loc_sram_buff_w14[15][4]}} & loc_sram_buff_w14[15][3:0]) | ({4{loc_sram_buff_w15[15][4]}} & loc_sram_buff_w15[15][3:0]);
	loc_rdata_buff[ 959: 956] = ({4{loc_sram_buff_w0[16][4]}} & loc_sram_buff_w0[16][3:0]) | ({4{loc_sram_buff_w1[16][4]}} & loc_sram_buff_w1[16][3:0]) | ({4{loc_sram_buff_w2[16][4]}} & loc_sram_buff_w2[16][3:0]) | ({4{loc_sram_buff_w3[16][4]}} & loc_sram_buff_w3[16][3:0]) | ({4{loc_sram_buff_w4[16][4]}} & loc_sram_buff_w4[16][3:0]) | ({4{loc_sram_buff_w5[16][4]}} & loc_sram_buff_w5[16][3:0]) | ({4{loc_sram_buff_w6[16][4]}} & loc_sram_buff_w6[16][3:0]) | ({4{loc_sram_buff_w7[16][4]}} & loc_sram_buff_w7[16][3:0]) | ({4{loc_sram_buff_w8[16][4]}} & loc_sram_buff_w8[16][3:0]) | ({4{loc_sram_buff_w9[16][4]}} & loc_sram_buff_w9[16][3:0]) | ({4{loc_sram_buff_w10[16][4]}} & loc_sram_buff_w10[16][3:0]) | ({4{loc_sram_buff_w11[16][4]}} & loc_sram_buff_w11[16][3:0]) | ({4{loc_sram_buff_w12[16][4]}} & loc_sram_buff_w12[16][3:0]) | ({4{loc_sram_buff_w13[16][4]}} & loc_sram_buff_w13[16][3:0]) | ({4{loc_sram_buff_w14[16][4]}} & loc_sram_buff_w14[16][3:0]) | ({4{loc_sram_buff_w15[16][4]}} & loc_sram_buff_w15[16][3:0]);
	loc_rdata_buff[ 955: 952] = ({4{loc_sram_buff_w0[17][4]}} & loc_sram_buff_w0[17][3:0]) | ({4{loc_sram_buff_w1[17][4]}} & loc_sram_buff_w1[17][3:0]) | ({4{loc_sram_buff_w2[17][4]}} & loc_sram_buff_w2[17][3:0]) | ({4{loc_sram_buff_w3[17][4]}} & loc_sram_buff_w3[17][3:0]) | ({4{loc_sram_buff_w4[17][4]}} & loc_sram_buff_w4[17][3:0]) | ({4{loc_sram_buff_w5[17][4]}} & loc_sram_buff_w5[17][3:0]) | ({4{loc_sram_buff_w6[17][4]}} & loc_sram_buff_w6[17][3:0]) | ({4{loc_sram_buff_w7[17][4]}} & loc_sram_buff_w7[17][3:0]) | ({4{loc_sram_buff_w8[17][4]}} & loc_sram_buff_w8[17][3:0]) | ({4{loc_sram_buff_w9[17][4]}} & loc_sram_buff_w9[17][3:0]) | ({4{loc_sram_buff_w10[17][4]}} & loc_sram_buff_w10[17][3:0]) | ({4{loc_sram_buff_w11[17][4]}} & loc_sram_buff_w11[17][3:0]) | ({4{loc_sram_buff_w12[17][4]}} & loc_sram_buff_w12[17][3:0]) | ({4{loc_sram_buff_w13[17][4]}} & loc_sram_buff_w13[17][3:0]) | ({4{loc_sram_buff_w14[17][4]}} & loc_sram_buff_w14[17][3:0]) | ({4{loc_sram_buff_w15[17][4]}} & loc_sram_buff_w15[17][3:0]);
	loc_rdata_buff[ 951: 948] = ({4{loc_sram_buff_w0[18][4]}} & loc_sram_buff_w0[18][3:0]) | ({4{loc_sram_buff_w1[18][4]}} & loc_sram_buff_w1[18][3:0]) | ({4{loc_sram_buff_w2[18][4]}} & loc_sram_buff_w2[18][3:0]) | ({4{loc_sram_buff_w3[18][4]}} & loc_sram_buff_w3[18][3:0]) | ({4{loc_sram_buff_w4[18][4]}} & loc_sram_buff_w4[18][3:0]) | ({4{loc_sram_buff_w5[18][4]}} & loc_sram_buff_w5[18][3:0]) | ({4{loc_sram_buff_w6[18][4]}} & loc_sram_buff_w6[18][3:0]) | ({4{loc_sram_buff_w7[18][4]}} & loc_sram_buff_w7[18][3:0]) | ({4{loc_sram_buff_w8[18][4]}} & loc_sram_buff_w8[18][3:0]) | ({4{loc_sram_buff_w9[18][4]}} & loc_sram_buff_w9[18][3:0]) | ({4{loc_sram_buff_w10[18][4]}} & loc_sram_buff_w10[18][3:0]) | ({4{loc_sram_buff_w11[18][4]}} & loc_sram_buff_w11[18][3:0]) | ({4{loc_sram_buff_w12[18][4]}} & loc_sram_buff_w12[18][3:0]) | ({4{loc_sram_buff_w13[18][4]}} & loc_sram_buff_w13[18][3:0]) | ({4{loc_sram_buff_w14[18][4]}} & loc_sram_buff_w14[18][3:0]) | ({4{loc_sram_buff_w15[18][4]}} & loc_sram_buff_w15[18][3:0]);
	loc_rdata_buff[ 947: 944] = ({4{loc_sram_buff_w0[19][4]}} & loc_sram_buff_w0[19][3:0]) | ({4{loc_sram_buff_w1[19][4]}} & loc_sram_buff_w1[19][3:0]) | ({4{loc_sram_buff_w2[19][4]}} & loc_sram_buff_w2[19][3:0]) | ({4{loc_sram_buff_w3[19][4]}} & loc_sram_buff_w3[19][3:0]) | ({4{loc_sram_buff_w4[19][4]}} & loc_sram_buff_w4[19][3:0]) | ({4{loc_sram_buff_w5[19][4]}} & loc_sram_buff_w5[19][3:0]) | ({4{loc_sram_buff_w6[19][4]}} & loc_sram_buff_w6[19][3:0]) | ({4{loc_sram_buff_w7[19][4]}} & loc_sram_buff_w7[19][3:0]) | ({4{loc_sram_buff_w8[19][4]}} & loc_sram_buff_w8[19][3:0]) | ({4{loc_sram_buff_w9[19][4]}} & loc_sram_buff_w9[19][3:0]) | ({4{loc_sram_buff_w10[19][4]}} & loc_sram_buff_w10[19][3:0]) | ({4{loc_sram_buff_w11[19][4]}} & loc_sram_buff_w11[19][3:0]) | ({4{loc_sram_buff_w12[19][4]}} & loc_sram_buff_w12[19][3:0]) | ({4{loc_sram_buff_w13[19][4]}} & loc_sram_buff_w13[19][3:0]) | ({4{loc_sram_buff_w14[19][4]}} & loc_sram_buff_w14[19][3:0]) | ({4{loc_sram_buff_w15[19][4]}} & loc_sram_buff_w15[19][3:0]);
	loc_rdata_buff[ 943: 940] = ({4{loc_sram_buff_w0[20][4]}} & loc_sram_buff_w0[20][3:0]) | ({4{loc_sram_buff_w1[20][4]}} & loc_sram_buff_w1[20][3:0]) | ({4{loc_sram_buff_w2[20][4]}} & loc_sram_buff_w2[20][3:0]) | ({4{loc_sram_buff_w3[20][4]}} & loc_sram_buff_w3[20][3:0]) | ({4{loc_sram_buff_w4[20][4]}} & loc_sram_buff_w4[20][3:0]) | ({4{loc_sram_buff_w5[20][4]}} & loc_sram_buff_w5[20][3:0]) | ({4{loc_sram_buff_w6[20][4]}} & loc_sram_buff_w6[20][3:0]) | ({4{loc_sram_buff_w7[20][4]}} & loc_sram_buff_w7[20][3:0]) | ({4{loc_sram_buff_w8[20][4]}} & loc_sram_buff_w8[20][3:0]) | ({4{loc_sram_buff_w9[20][4]}} & loc_sram_buff_w9[20][3:0]) | ({4{loc_sram_buff_w10[20][4]}} & loc_sram_buff_w10[20][3:0]) | ({4{loc_sram_buff_w11[20][4]}} & loc_sram_buff_w11[20][3:0]) | ({4{loc_sram_buff_w12[20][4]}} & loc_sram_buff_w12[20][3:0]) | ({4{loc_sram_buff_w13[20][4]}} & loc_sram_buff_w13[20][3:0]) | ({4{loc_sram_buff_w14[20][4]}} & loc_sram_buff_w14[20][3:0]) | ({4{loc_sram_buff_w15[20][4]}} & loc_sram_buff_w15[20][3:0]);
	loc_rdata_buff[ 939: 936] = ({4{loc_sram_buff_w0[21][4]}} & loc_sram_buff_w0[21][3:0]) | ({4{loc_sram_buff_w1[21][4]}} & loc_sram_buff_w1[21][3:0]) | ({4{loc_sram_buff_w2[21][4]}} & loc_sram_buff_w2[21][3:0]) | ({4{loc_sram_buff_w3[21][4]}} & loc_sram_buff_w3[21][3:0]) | ({4{loc_sram_buff_w4[21][4]}} & loc_sram_buff_w4[21][3:0]) | ({4{loc_sram_buff_w5[21][4]}} & loc_sram_buff_w5[21][3:0]) | ({4{loc_sram_buff_w6[21][4]}} & loc_sram_buff_w6[21][3:0]) | ({4{loc_sram_buff_w7[21][4]}} & loc_sram_buff_w7[21][3:0]) | ({4{loc_sram_buff_w8[21][4]}} & loc_sram_buff_w8[21][3:0]) | ({4{loc_sram_buff_w9[21][4]}} & loc_sram_buff_w9[21][3:0]) | ({4{loc_sram_buff_w10[21][4]}} & loc_sram_buff_w10[21][3:0]) | ({4{loc_sram_buff_w11[21][4]}} & loc_sram_buff_w11[21][3:0]) | ({4{loc_sram_buff_w12[21][4]}} & loc_sram_buff_w12[21][3:0]) | ({4{loc_sram_buff_w13[21][4]}} & loc_sram_buff_w13[21][3:0]) | ({4{loc_sram_buff_w14[21][4]}} & loc_sram_buff_w14[21][3:0]) | ({4{loc_sram_buff_w15[21][4]}} & loc_sram_buff_w15[21][3:0]);
	loc_rdata_buff[ 935: 932] = ({4{loc_sram_buff_w0[22][4]}} & loc_sram_buff_w0[22][3:0]) | ({4{loc_sram_buff_w1[22][4]}} & loc_sram_buff_w1[22][3:0]) | ({4{loc_sram_buff_w2[22][4]}} & loc_sram_buff_w2[22][3:0]) | ({4{loc_sram_buff_w3[22][4]}} & loc_sram_buff_w3[22][3:0]) | ({4{loc_sram_buff_w4[22][4]}} & loc_sram_buff_w4[22][3:0]) | ({4{loc_sram_buff_w5[22][4]}} & loc_sram_buff_w5[22][3:0]) | ({4{loc_sram_buff_w6[22][4]}} & loc_sram_buff_w6[22][3:0]) | ({4{loc_sram_buff_w7[22][4]}} & loc_sram_buff_w7[22][3:0]) | ({4{loc_sram_buff_w8[22][4]}} & loc_sram_buff_w8[22][3:0]) | ({4{loc_sram_buff_w9[22][4]}} & loc_sram_buff_w9[22][3:0]) | ({4{loc_sram_buff_w10[22][4]}} & loc_sram_buff_w10[22][3:0]) | ({4{loc_sram_buff_w11[22][4]}} & loc_sram_buff_w11[22][3:0]) | ({4{loc_sram_buff_w12[22][4]}} & loc_sram_buff_w12[22][3:0]) | ({4{loc_sram_buff_w13[22][4]}} & loc_sram_buff_w13[22][3:0]) | ({4{loc_sram_buff_w14[22][4]}} & loc_sram_buff_w14[22][3:0]) | ({4{loc_sram_buff_w15[22][4]}} & loc_sram_buff_w15[22][3:0]);
	loc_rdata_buff[ 931: 928] = ({4{loc_sram_buff_w0[23][4]}} & loc_sram_buff_w0[23][3:0]) | ({4{loc_sram_buff_w1[23][4]}} & loc_sram_buff_w1[23][3:0]) | ({4{loc_sram_buff_w2[23][4]}} & loc_sram_buff_w2[23][3:0]) | ({4{loc_sram_buff_w3[23][4]}} & loc_sram_buff_w3[23][3:0]) | ({4{loc_sram_buff_w4[23][4]}} & loc_sram_buff_w4[23][3:0]) | ({4{loc_sram_buff_w5[23][4]}} & loc_sram_buff_w5[23][3:0]) | ({4{loc_sram_buff_w6[23][4]}} & loc_sram_buff_w6[23][3:0]) | ({4{loc_sram_buff_w7[23][4]}} & loc_sram_buff_w7[23][3:0]) | ({4{loc_sram_buff_w8[23][4]}} & loc_sram_buff_w8[23][3:0]) | ({4{loc_sram_buff_w9[23][4]}} & loc_sram_buff_w9[23][3:0]) | ({4{loc_sram_buff_w10[23][4]}} & loc_sram_buff_w10[23][3:0]) | ({4{loc_sram_buff_w11[23][4]}} & loc_sram_buff_w11[23][3:0]) | ({4{loc_sram_buff_w12[23][4]}} & loc_sram_buff_w12[23][3:0]) | ({4{loc_sram_buff_w13[23][4]}} & loc_sram_buff_w13[23][3:0]) | ({4{loc_sram_buff_w14[23][4]}} & loc_sram_buff_w14[23][3:0]) | ({4{loc_sram_buff_w15[23][4]}} & loc_sram_buff_w15[23][3:0]);
	loc_rdata_buff[ 927: 924] = ({4{loc_sram_buff_w0[24][4]}} & loc_sram_buff_w0[24][3:0]) | ({4{loc_sram_buff_w1[24][4]}} & loc_sram_buff_w1[24][3:0]) | ({4{loc_sram_buff_w2[24][4]}} & loc_sram_buff_w2[24][3:0]) | ({4{loc_sram_buff_w3[24][4]}} & loc_sram_buff_w3[24][3:0]) | ({4{loc_sram_buff_w4[24][4]}} & loc_sram_buff_w4[24][3:0]) | ({4{loc_sram_buff_w5[24][4]}} & loc_sram_buff_w5[24][3:0]) | ({4{loc_sram_buff_w6[24][4]}} & loc_sram_buff_w6[24][3:0]) | ({4{loc_sram_buff_w7[24][4]}} & loc_sram_buff_w7[24][3:0]) | ({4{loc_sram_buff_w8[24][4]}} & loc_sram_buff_w8[24][3:0]) | ({4{loc_sram_buff_w9[24][4]}} & loc_sram_buff_w9[24][3:0]) | ({4{loc_sram_buff_w10[24][4]}} & loc_sram_buff_w10[24][3:0]) | ({4{loc_sram_buff_w11[24][4]}} & loc_sram_buff_w11[24][3:0]) | ({4{loc_sram_buff_w12[24][4]}} & loc_sram_buff_w12[24][3:0]) | ({4{loc_sram_buff_w13[24][4]}} & loc_sram_buff_w13[24][3:0]) | ({4{loc_sram_buff_w14[24][4]}} & loc_sram_buff_w14[24][3:0]) | ({4{loc_sram_buff_w15[24][4]}} & loc_sram_buff_w15[24][3:0]);
	loc_rdata_buff[ 923: 920] = ({4{loc_sram_buff_w0[25][4]}} & loc_sram_buff_w0[25][3:0]) | ({4{loc_sram_buff_w1[25][4]}} & loc_sram_buff_w1[25][3:0]) | ({4{loc_sram_buff_w2[25][4]}} & loc_sram_buff_w2[25][3:0]) | ({4{loc_sram_buff_w3[25][4]}} & loc_sram_buff_w3[25][3:0]) | ({4{loc_sram_buff_w4[25][4]}} & loc_sram_buff_w4[25][3:0]) | ({4{loc_sram_buff_w5[25][4]}} & loc_sram_buff_w5[25][3:0]) | ({4{loc_sram_buff_w6[25][4]}} & loc_sram_buff_w6[25][3:0]) | ({4{loc_sram_buff_w7[25][4]}} & loc_sram_buff_w7[25][3:0]) | ({4{loc_sram_buff_w8[25][4]}} & loc_sram_buff_w8[25][3:0]) | ({4{loc_sram_buff_w9[25][4]}} & loc_sram_buff_w9[25][3:0]) | ({4{loc_sram_buff_w10[25][4]}} & loc_sram_buff_w10[25][3:0]) | ({4{loc_sram_buff_w11[25][4]}} & loc_sram_buff_w11[25][3:0]) | ({4{loc_sram_buff_w12[25][4]}} & loc_sram_buff_w12[25][3:0]) | ({4{loc_sram_buff_w13[25][4]}} & loc_sram_buff_w13[25][3:0]) | ({4{loc_sram_buff_w14[25][4]}} & loc_sram_buff_w14[25][3:0]) | ({4{loc_sram_buff_w15[25][4]}} & loc_sram_buff_w15[25][3:0]);
	loc_rdata_buff[ 919: 916] = ({4{loc_sram_buff_w0[26][4]}} & loc_sram_buff_w0[26][3:0]) | ({4{loc_sram_buff_w1[26][4]}} & loc_sram_buff_w1[26][3:0]) | ({4{loc_sram_buff_w2[26][4]}} & loc_sram_buff_w2[26][3:0]) | ({4{loc_sram_buff_w3[26][4]}} & loc_sram_buff_w3[26][3:0]) | ({4{loc_sram_buff_w4[26][4]}} & loc_sram_buff_w4[26][3:0]) | ({4{loc_sram_buff_w5[26][4]}} & loc_sram_buff_w5[26][3:0]) | ({4{loc_sram_buff_w6[26][4]}} & loc_sram_buff_w6[26][3:0]) | ({4{loc_sram_buff_w7[26][4]}} & loc_sram_buff_w7[26][3:0]) | ({4{loc_sram_buff_w8[26][4]}} & loc_sram_buff_w8[26][3:0]) | ({4{loc_sram_buff_w9[26][4]}} & loc_sram_buff_w9[26][3:0]) | ({4{loc_sram_buff_w10[26][4]}} & loc_sram_buff_w10[26][3:0]) | ({4{loc_sram_buff_w11[26][4]}} & loc_sram_buff_w11[26][3:0]) | ({4{loc_sram_buff_w12[26][4]}} & loc_sram_buff_w12[26][3:0]) | ({4{loc_sram_buff_w13[26][4]}} & loc_sram_buff_w13[26][3:0]) | ({4{loc_sram_buff_w14[26][4]}} & loc_sram_buff_w14[26][3:0]) | ({4{loc_sram_buff_w15[26][4]}} & loc_sram_buff_w15[26][3:0]);
	loc_rdata_buff[ 915: 912] = ({4{loc_sram_buff_w0[27][4]}} & loc_sram_buff_w0[27][3:0]) | ({4{loc_sram_buff_w1[27][4]}} & loc_sram_buff_w1[27][3:0]) | ({4{loc_sram_buff_w2[27][4]}} & loc_sram_buff_w2[27][3:0]) | ({4{loc_sram_buff_w3[27][4]}} & loc_sram_buff_w3[27][3:0]) | ({4{loc_sram_buff_w4[27][4]}} & loc_sram_buff_w4[27][3:0]) | ({4{loc_sram_buff_w5[27][4]}} & loc_sram_buff_w5[27][3:0]) | ({4{loc_sram_buff_w6[27][4]}} & loc_sram_buff_w6[27][3:0]) | ({4{loc_sram_buff_w7[27][4]}} & loc_sram_buff_w7[27][3:0]) | ({4{loc_sram_buff_w8[27][4]}} & loc_sram_buff_w8[27][3:0]) | ({4{loc_sram_buff_w9[27][4]}} & loc_sram_buff_w9[27][3:0]) | ({4{loc_sram_buff_w10[27][4]}} & loc_sram_buff_w10[27][3:0]) | ({4{loc_sram_buff_w11[27][4]}} & loc_sram_buff_w11[27][3:0]) | ({4{loc_sram_buff_w12[27][4]}} & loc_sram_buff_w12[27][3:0]) | ({4{loc_sram_buff_w13[27][4]}} & loc_sram_buff_w13[27][3:0]) | ({4{loc_sram_buff_w14[27][4]}} & loc_sram_buff_w14[27][3:0]) | ({4{loc_sram_buff_w15[27][4]}} & loc_sram_buff_w15[27][3:0]);
	loc_rdata_buff[ 911: 908] = ({4{loc_sram_buff_w0[28][4]}} & loc_sram_buff_w0[28][3:0]) | ({4{loc_sram_buff_w1[28][4]}} & loc_sram_buff_w1[28][3:0]) | ({4{loc_sram_buff_w2[28][4]}} & loc_sram_buff_w2[28][3:0]) | ({4{loc_sram_buff_w3[28][4]}} & loc_sram_buff_w3[28][3:0]) | ({4{loc_sram_buff_w4[28][4]}} & loc_sram_buff_w4[28][3:0]) | ({4{loc_sram_buff_w5[28][4]}} & loc_sram_buff_w5[28][3:0]) | ({4{loc_sram_buff_w6[28][4]}} & loc_sram_buff_w6[28][3:0]) | ({4{loc_sram_buff_w7[28][4]}} & loc_sram_buff_w7[28][3:0]) | ({4{loc_sram_buff_w8[28][4]}} & loc_sram_buff_w8[28][3:0]) | ({4{loc_sram_buff_w9[28][4]}} & loc_sram_buff_w9[28][3:0]) | ({4{loc_sram_buff_w10[28][4]}} & loc_sram_buff_w10[28][3:0]) | ({4{loc_sram_buff_w11[28][4]}} & loc_sram_buff_w11[28][3:0]) | ({4{loc_sram_buff_w12[28][4]}} & loc_sram_buff_w12[28][3:0]) | ({4{loc_sram_buff_w13[28][4]}} & loc_sram_buff_w13[28][3:0]) | ({4{loc_sram_buff_w14[28][4]}} & loc_sram_buff_w14[28][3:0]) | ({4{loc_sram_buff_w15[28][4]}} & loc_sram_buff_w15[28][3:0]);
	loc_rdata_buff[ 907: 904] = ({4{loc_sram_buff_w0[29][4]}} & loc_sram_buff_w0[29][3:0]) | ({4{loc_sram_buff_w1[29][4]}} & loc_sram_buff_w1[29][3:0]) | ({4{loc_sram_buff_w2[29][4]}} & loc_sram_buff_w2[29][3:0]) | ({4{loc_sram_buff_w3[29][4]}} & loc_sram_buff_w3[29][3:0]) | ({4{loc_sram_buff_w4[29][4]}} & loc_sram_buff_w4[29][3:0]) | ({4{loc_sram_buff_w5[29][4]}} & loc_sram_buff_w5[29][3:0]) | ({4{loc_sram_buff_w6[29][4]}} & loc_sram_buff_w6[29][3:0]) | ({4{loc_sram_buff_w7[29][4]}} & loc_sram_buff_w7[29][3:0]) | ({4{loc_sram_buff_w8[29][4]}} & loc_sram_buff_w8[29][3:0]) | ({4{loc_sram_buff_w9[29][4]}} & loc_sram_buff_w9[29][3:0]) | ({4{loc_sram_buff_w10[29][4]}} & loc_sram_buff_w10[29][3:0]) | ({4{loc_sram_buff_w11[29][4]}} & loc_sram_buff_w11[29][3:0]) | ({4{loc_sram_buff_w12[29][4]}} & loc_sram_buff_w12[29][3:0]) | ({4{loc_sram_buff_w13[29][4]}} & loc_sram_buff_w13[29][3:0]) | ({4{loc_sram_buff_w14[29][4]}} & loc_sram_buff_w14[29][3:0]) | ({4{loc_sram_buff_w15[29][4]}} & loc_sram_buff_w15[29][3:0]);
	loc_rdata_buff[ 903: 900] = ({4{loc_sram_buff_w0[30][4]}} & loc_sram_buff_w0[30][3:0]) | ({4{loc_sram_buff_w1[30][4]}} & loc_sram_buff_w1[30][3:0]) | ({4{loc_sram_buff_w2[30][4]}} & loc_sram_buff_w2[30][3:0]) | ({4{loc_sram_buff_w3[30][4]}} & loc_sram_buff_w3[30][3:0]) | ({4{loc_sram_buff_w4[30][4]}} & loc_sram_buff_w4[30][3:0]) | ({4{loc_sram_buff_w5[30][4]}} & loc_sram_buff_w5[30][3:0]) | ({4{loc_sram_buff_w6[30][4]}} & loc_sram_buff_w6[30][3:0]) | ({4{loc_sram_buff_w7[30][4]}} & loc_sram_buff_w7[30][3:0]) | ({4{loc_sram_buff_w8[30][4]}} & loc_sram_buff_w8[30][3:0]) | ({4{loc_sram_buff_w9[30][4]}} & loc_sram_buff_w9[30][3:0]) | ({4{loc_sram_buff_w10[30][4]}} & loc_sram_buff_w10[30][3:0]) | ({4{loc_sram_buff_w11[30][4]}} & loc_sram_buff_w11[30][3:0]) | ({4{loc_sram_buff_w12[30][4]}} & loc_sram_buff_w12[30][3:0]) | ({4{loc_sram_buff_w13[30][4]}} & loc_sram_buff_w13[30][3:0]) | ({4{loc_sram_buff_w14[30][4]}} & loc_sram_buff_w14[30][3:0]) | ({4{loc_sram_buff_w15[30][4]}} & loc_sram_buff_w15[30][3:0]);
	loc_rdata_buff[ 899: 896] = ({4{loc_sram_buff_w0[31][4]}} & loc_sram_buff_w0[31][3:0]) | ({4{loc_sram_buff_w1[31][4]}} & loc_sram_buff_w1[31][3:0]) | ({4{loc_sram_buff_w2[31][4]}} & loc_sram_buff_w2[31][3:0]) | ({4{loc_sram_buff_w3[31][4]}} & loc_sram_buff_w3[31][3:0]) | ({4{loc_sram_buff_w4[31][4]}} & loc_sram_buff_w4[31][3:0]) | ({4{loc_sram_buff_w5[31][4]}} & loc_sram_buff_w5[31][3:0]) | ({4{loc_sram_buff_w6[31][4]}} & loc_sram_buff_w6[31][3:0]) | ({4{loc_sram_buff_w7[31][4]}} & loc_sram_buff_w7[31][3:0]) | ({4{loc_sram_buff_w8[31][4]}} & loc_sram_buff_w8[31][3:0]) | ({4{loc_sram_buff_w9[31][4]}} & loc_sram_buff_w9[31][3:0]) | ({4{loc_sram_buff_w10[31][4]}} & loc_sram_buff_w10[31][3:0]) | ({4{loc_sram_buff_w11[31][4]}} & loc_sram_buff_w11[31][3:0]) | ({4{loc_sram_buff_w12[31][4]}} & loc_sram_buff_w12[31][3:0]) | ({4{loc_sram_buff_w13[31][4]}} & loc_sram_buff_w13[31][3:0]) | ({4{loc_sram_buff_w14[31][4]}} & loc_sram_buff_w14[31][3:0]) | ({4{loc_sram_buff_w15[31][4]}} & loc_sram_buff_w15[31][3:0]);
	loc_rdata_buff[ 895: 892] = ({4{loc_sram_buff_w0[32][4]}} & loc_sram_buff_w0[32][3:0]) | ({4{loc_sram_buff_w1[32][4]}} & loc_sram_buff_w1[32][3:0]) | ({4{loc_sram_buff_w2[32][4]}} & loc_sram_buff_w2[32][3:0]) | ({4{loc_sram_buff_w3[32][4]}} & loc_sram_buff_w3[32][3:0]) | ({4{loc_sram_buff_w4[32][4]}} & loc_sram_buff_w4[32][3:0]) | ({4{loc_sram_buff_w5[32][4]}} & loc_sram_buff_w5[32][3:0]) | ({4{loc_sram_buff_w6[32][4]}} & loc_sram_buff_w6[32][3:0]) | ({4{loc_sram_buff_w7[32][4]}} & loc_sram_buff_w7[32][3:0]) | ({4{loc_sram_buff_w8[32][4]}} & loc_sram_buff_w8[32][3:0]) | ({4{loc_sram_buff_w9[32][4]}} & loc_sram_buff_w9[32][3:0]) | ({4{loc_sram_buff_w10[32][4]}} & loc_sram_buff_w10[32][3:0]) | ({4{loc_sram_buff_w11[32][4]}} & loc_sram_buff_w11[32][3:0]) | ({4{loc_sram_buff_w12[32][4]}} & loc_sram_buff_w12[32][3:0]) | ({4{loc_sram_buff_w13[32][4]}} & loc_sram_buff_w13[32][3:0]) | ({4{loc_sram_buff_w14[32][4]}} & loc_sram_buff_w14[32][3:0]) | ({4{loc_sram_buff_w15[32][4]}} & loc_sram_buff_w15[32][3:0]);
	loc_rdata_buff[ 891: 888] = ({4{loc_sram_buff_w0[33][4]}} & loc_sram_buff_w0[33][3:0]) | ({4{loc_sram_buff_w1[33][4]}} & loc_sram_buff_w1[33][3:0]) | ({4{loc_sram_buff_w2[33][4]}} & loc_sram_buff_w2[33][3:0]) | ({4{loc_sram_buff_w3[33][4]}} & loc_sram_buff_w3[33][3:0]) | ({4{loc_sram_buff_w4[33][4]}} & loc_sram_buff_w4[33][3:0]) | ({4{loc_sram_buff_w5[33][4]}} & loc_sram_buff_w5[33][3:0]) | ({4{loc_sram_buff_w6[33][4]}} & loc_sram_buff_w6[33][3:0]) | ({4{loc_sram_buff_w7[33][4]}} & loc_sram_buff_w7[33][3:0]) | ({4{loc_sram_buff_w8[33][4]}} & loc_sram_buff_w8[33][3:0]) | ({4{loc_sram_buff_w9[33][4]}} & loc_sram_buff_w9[33][3:0]) | ({4{loc_sram_buff_w10[33][4]}} & loc_sram_buff_w10[33][3:0]) | ({4{loc_sram_buff_w11[33][4]}} & loc_sram_buff_w11[33][3:0]) | ({4{loc_sram_buff_w12[33][4]}} & loc_sram_buff_w12[33][3:0]) | ({4{loc_sram_buff_w13[33][4]}} & loc_sram_buff_w13[33][3:0]) | ({4{loc_sram_buff_w14[33][4]}} & loc_sram_buff_w14[33][3:0]) | ({4{loc_sram_buff_w15[33][4]}} & loc_sram_buff_w15[33][3:0]);
	loc_rdata_buff[ 887: 884] = ({4{loc_sram_buff_w0[34][4]}} & loc_sram_buff_w0[34][3:0]) | ({4{loc_sram_buff_w1[34][4]}} & loc_sram_buff_w1[34][3:0]) | ({4{loc_sram_buff_w2[34][4]}} & loc_sram_buff_w2[34][3:0]) | ({4{loc_sram_buff_w3[34][4]}} & loc_sram_buff_w3[34][3:0]) | ({4{loc_sram_buff_w4[34][4]}} & loc_sram_buff_w4[34][3:0]) | ({4{loc_sram_buff_w5[34][4]}} & loc_sram_buff_w5[34][3:0]) | ({4{loc_sram_buff_w6[34][4]}} & loc_sram_buff_w6[34][3:0]) | ({4{loc_sram_buff_w7[34][4]}} & loc_sram_buff_w7[34][3:0]) | ({4{loc_sram_buff_w8[34][4]}} & loc_sram_buff_w8[34][3:0]) | ({4{loc_sram_buff_w9[34][4]}} & loc_sram_buff_w9[34][3:0]) | ({4{loc_sram_buff_w10[34][4]}} & loc_sram_buff_w10[34][3:0]) | ({4{loc_sram_buff_w11[34][4]}} & loc_sram_buff_w11[34][3:0]) | ({4{loc_sram_buff_w12[34][4]}} & loc_sram_buff_w12[34][3:0]) | ({4{loc_sram_buff_w13[34][4]}} & loc_sram_buff_w13[34][3:0]) | ({4{loc_sram_buff_w14[34][4]}} & loc_sram_buff_w14[34][3:0]) | ({4{loc_sram_buff_w15[34][4]}} & loc_sram_buff_w15[34][3:0]);
	loc_rdata_buff[ 883: 880] = ({4{loc_sram_buff_w0[35][4]}} & loc_sram_buff_w0[35][3:0]) | ({4{loc_sram_buff_w1[35][4]}} & loc_sram_buff_w1[35][3:0]) | ({4{loc_sram_buff_w2[35][4]}} & loc_sram_buff_w2[35][3:0]) | ({4{loc_sram_buff_w3[35][4]}} & loc_sram_buff_w3[35][3:0]) | ({4{loc_sram_buff_w4[35][4]}} & loc_sram_buff_w4[35][3:0]) | ({4{loc_sram_buff_w5[35][4]}} & loc_sram_buff_w5[35][3:0]) | ({4{loc_sram_buff_w6[35][4]}} & loc_sram_buff_w6[35][3:0]) | ({4{loc_sram_buff_w7[35][4]}} & loc_sram_buff_w7[35][3:0]) | ({4{loc_sram_buff_w8[35][4]}} & loc_sram_buff_w8[35][3:0]) | ({4{loc_sram_buff_w9[35][4]}} & loc_sram_buff_w9[35][3:0]) | ({4{loc_sram_buff_w10[35][4]}} & loc_sram_buff_w10[35][3:0]) | ({4{loc_sram_buff_w11[35][4]}} & loc_sram_buff_w11[35][3:0]) | ({4{loc_sram_buff_w12[35][4]}} & loc_sram_buff_w12[35][3:0]) | ({4{loc_sram_buff_w13[35][4]}} & loc_sram_buff_w13[35][3:0]) | ({4{loc_sram_buff_w14[35][4]}} & loc_sram_buff_w14[35][3:0]) | ({4{loc_sram_buff_w15[35][4]}} & loc_sram_buff_w15[35][3:0]);
	loc_rdata_buff[ 879: 876] = ({4{loc_sram_buff_w0[36][4]}} & loc_sram_buff_w0[36][3:0]) | ({4{loc_sram_buff_w1[36][4]}} & loc_sram_buff_w1[36][3:0]) | ({4{loc_sram_buff_w2[36][4]}} & loc_sram_buff_w2[36][3:0]) | ({4{loc_sram_buff_w3[36][4]}} & loc_sram_buff_w3[36][3:0]) | ({4{loc_sram_buff_w4[36][4]}} & loc_sram_buff_w4[36][3:0]) | ({4{loc_sram_buff_w5[36][4]}} & loc_sram_buff_w5[36][3:0]) | ({4{loc_sram_buff_w6[36][4]}} & loc_sram_buff_w6[36][3:0]) | ({4{loc_sram_buff_w7[36][4]}} & loc_sram_buff_w7[36][3:0]) | ({4{loc_sram_buff_w8[36][4]}} & loc_sram_buff_w8[36][3:0]) | ({4{loc_sram_buff_w9[36][4]}} & loc_sram_buff_w9[36][3:0]) | ({4{loc_sram_buff_w10[36][4]}} & loc_sram_buff_w10[36][3:0]) | ({4{loc_sram_buff_w11[36][4]}} & loc_sram_buff_w11[36][3:0]) | ({4{loc_sram_buff_w12[36][4]}} & loc_sram_buff_w12[36][3:0]) | ({4{loc_sram_buff_w13[36][4]}} & loc_sram_buff_w13[36][3:0]) | ({4{loc_sram_buff_w14[36][4]}} & loc_sram_buff_w14[36][3:0]) | ({4{loc_sram_buff_w15[36][4]}} & loc_sram_buff_w15[36][3:0]);
	loc_rdata_buff[ 875: 872] = ({4{loc_sram_buff_w0[37][4]}} & loc_sram_buff_w0[37][3:0]) | ({4{loc_sram_buff_w1[37][4]}} & loc_sram_buff_w1[37][3:0]) | ({4{loc_sram_buff_w2[37][4]}} & loc_sram_buff_w2[37][3:0]) | ({4{loc_sram_buff_w3[37][4]}} & loc_sram_buff_w3[37][3:0]) | ({4{loc_sram_buff_w4[37][4]}} & loc_sram_buff_w4[37][3:0]) | ({4{loc_sram_buff_w5[37][4]}} & loc_sram_buff_w5[37][3:0]) | ({4{loc_sram_buff_w6[37][4]}} & loc_sram_buff_w6[37][3:0]) | ({4{loc_sram_buff_w7[37][4]}} & loc_sram_buff_w7[37][3:0]) | ({4{loc_sram_buff_w8[37][4]}} & loc_sram_buff_w8[37][3:0]) | ({4{loc_sram_buff_w9[37][4]}} & loc_sram_buff_w9[37][3:0]) | ({4{loc_sram_buff_w10[37][4]}} & loc_sram_buff_w10[37][3:0]) | ({4{loc_sram_buff_w11[37][4]}} & loc_sram_buff_w11[37][3:0]) | ({4{loc_sram_buff_w12[37][4]}} & loc_sram_buff_w12[37][3:0]) | ({4{loc_sram_buff_w13[37][4]}} & loc_sram_buff_w13[37][3:0]) | ({4{loc_sram_buff_w14[37][4]}} & loc_sram_buff_w14[37][3:0]) | ({4{loc_sram_buff_w15[37][4]}} & loc_sram_buff_w15[37][3:0]);
	loc_rdata_buff[ 871: 868] = ({4{loc_sram_buff_w0[38][4]}} & loc_sram_buff_w0[38][3:0]) | ({4{loc_sram_buff_w1[38][4]}} & loc_sram_buff_w1[38][3:0]) | ({4{loc_sram_buff_w2[38][4]}} & loc_sram_buff_w2[38][3:0]) | ({4{loc_sram_buff_w3[38][4]}} & loc_sram_buff_w3[38][3:0]) | ({4{loc_sram_buff_w4[38][4]}} & loc_sram_buff_w4[38][3:0]) | ({4{loc_sram_buff_w5[38][4]}} & loc_sram_buff_w5[38][3:0]) | ({4{loc_sram_buff_w6[38][4]}} & loc_sram_buff_w6[38][3:0]) | ({4{loc_sram_buff_w7[38][4]}} & loc_sram_buff_w7[38][3:0]) | ({4{loc_sram_buff_w8[38][4]}} & loc_sram_buff_w8[38][3:0]) | ({4{loc_sram_buff_w9[38][4]}} & loc_sram_buff_w9[38][3:0]) | ({4{loc_sram_buff_w10[38][4]}} & loc_sram_buff_w10[38][3:0]) | ({4{loc_sram_buff_w11[38][4]}} & loc_sram_buff_w11[38][3:0]) | ({4{loc_sram_buff_w12[38][4]}} & loc_sram_buff_w12[38][3:0]) | ({4{loc_sram_buff_w13[38][4]}} & loc_sram_buff_w13[38][3:0]) | ({4{loc_sram_buff_w14[38][4]}} & loc_sram_buff_w14[38][3:0]) | ({4{loc_sram_buff_w15[38][4]}} & loc_sram_buff_w15[38][3:0]);
	loc_rdata_buff[ 867: 864] = ({4{loc_sram_buff_w0[39][4]}} & loc_sram_buff_w0[39][3:0]) | ({4{loc_sram_buff_w1[39][4]}} & loc_sram_buff_w1[39][3:0]) | ({4{loc_sram_buff_w2[39][4]}} & loc_sram_buff_w2[39][3:0]) | ({4{loc_sram_buff_w3[39][4]}} & loc_sram_buff_w3[39][3:0]) | ({4{loc_sram_buff_w4[39][4]}} & loc_sram_buff_w4[39][3:0]) | ({4{loc_sram_buff_w5[39][4]}} & loc_sram_buff_w5[39][3:0]) | ({4{loc_sram_buff_w6[39][4]}} & loc_sram_buff_w6[39][3:0]) | ({4{loc_sram_buff_w7[39][4]}} & loc_sram_buff_w7[39][3:0]) | ({4{loc_sram_buff_w8[39][4]}} & loc_sram_buff_w8[39][3:0]) | ({4{loc_sram_buff_w9[39][4]}} & loc_sram_buff_w9[39][3:0]) | ({4{loc_sram_buff_w10[39][4]}} & loc_sram_buff_w10[39][3:0]) | ({4{loc_sram_buff_w11[39][4]}} & loc_sram_buff_w11[39][3:0]) | ({4{loc_sram_buff_w12[39][4]}} & loc_sram_buff_w12[39][3:0]) | ({4{loc_sram_buff_w13[39][4]}} & loc_sram_buff_w13[39][3:0]) | ({4{loc_sram_buff_w14[39][4]}} & loc_sram_buff_w14[39][3:0]) | ({4{loc_sram_buff_w15[39][4]}} & loc_sram_buff_w15[39][3:0]);
	loc_rdata_buff[ 863: 860] = ({4{loc_sram_buff_w0[40][4]}} & loc_sram_buff_w0[40][3:0]) | ({4{loc_sram_buff_w1[40][4]}} & loc_sram_buff_w1[40][3:0]) | ({4{loc_sram_buff_w2[40][4]}} & loc_sram_buff_w2[40][3:0]) | ({4{loc_sram_buff_w3[40][4]}} & loc_sram_buff_w3[40][3:0]) | ({4{loc_sram_buff_w4[40][4]}} & loc_sram_buff_w4[40][3:0]) | ({4{loc_sram_buff_w5[40][4]}} & loc_sram_buff_w5[40][3:0]) | ({4{loc_sram_buff_w6[40][4]}} & loc_sram_buff_w6[40][3:0]) | ({4{loc_sram_buff_w7[40][4]}} & loc_sram_buff_w7[40][3:0]) | ({4{loc_sram_buff_w8[40][4]}} & loc_sram_buff_w8[40][3:0]) | ({4{loc_sram_buff_w9[40][4]}} & loc_sram_buff_w9[40][3:0]) | ({4{loc_sram_buff_w10[40][4]}} & loc_sram_buff_w10[40][3:0]) | ({4{loc_sram_buff_w11[40][4]}} & loc_sram_buff_w11[40][3:0]) | ({4{loc_sram_buff_w12[40][4]}} & loc_sram_buff_w12[40][3:0]) | ({4{loc_sram_buff_w13[40][4]}} & loc_sram_buff_w13[40][3:0]) | ({4{loc_sram_buff_w14[40][4]}} & loc_sram_buff_w14[40][3:0]) | ({4{loc_sram_buff_w15[40][4]}} & loc_sram_buff_w15[40][3:0]);
	loc_rdata_buff[ 859: 856] = ({4{loc_sram_buff_w0[41][4]}} & loc_sram_buff_w0[41][3:0]) | ({4{loc_sram_buff_w1[41][4]}} & loc_sram_buff_w1[41][3:0]) | ({4{loc_sram_buff_w2[41][4]}} & loc_sram_buff_w2[41][3:0]) | ({4{loc_sram_buff_w3[41][4]}} & loc_sram_buff_w3[41][3:0]) | ({4{loc_sram_buff_w4[41][4]}} & loc_sram_buff_w4[41][3:0]) | ({4{loc_sram_buff_w5[41][4]}} & loc_sram_buff_w5[41][3:0]) | ({4{loc_sram_buff_w6[41][4]}} & loc_sram_buff_w6[41][3:0]) | ({4{loc_sram_buff_w7[41][4]}} & loc_sram_buff_w7[41][3:0]) | ({4{loc_sram_buff_w8[41][4]}} & loc_sram_buff_w8[41][3:0]) | ({4{loc_sram_buff_w9[41][4]}} & loc_sram_buff_w9[41][3:0]) | ({4{loc_sram_buff_w10[41][4]}} & loc_sram_buff_w10[41][3:0]) | ({4{loc_sram_buff_w11[41][4]}} & loc_sram_buff_w11[41][3:0]) | ({4{loc_sram_buff_w12[41][4]}} & loc_sram_buff_w12[41][3:0]) | ({4{loc_sram_buff_w13[41][4]}} & loc_sram_buff_w13[41][3:0]) | ({4{loc_sram_buff_w14[41][4]}} & loc_sram_buff_w14[41][3:0]) | ({4{loc_sram_buff_w15[41][4]}} & loc_sram_buff_w15[41][3:0]);
	loc_rdata_buff[ 855: 852] = ({4{loc_sram_buff_w0[42][4]}} & loc_sram_buff_w0[42][3:0]) | ({4{loc_sram_buff_w1[42][4]}} & loc_sram_buff_w1[42][3:0]) | ({4{loc_sram_buff_w2[42][4]}} & loc_sram_buff_w2[42][3:0]) | ({4{loc_sram_buff_w3[42][4]}} & loc_sram_buff_w3[42][3:0]) | ({4{loc_sram_buff_w4[42][4]}} & loc_sram_buff_w4[42][3:0]) | ({4{loc_sram_buff_w5[42][4]}} & loc_sram_buff_w5[42][3:0]) | ({4{loc_sram_buff_w6[42][4]}} & loc_sram_buff_w6[42][3:0]) | ({4{loc_sram_buff_w7[42][4]}} & loc_sram_buff_w7[42][3:0]) | ({4{loc_sram_buff_w8[42][4]}} & loc_sram_buff_w8[42][3:0]) | ({4{loc_sram_buff_w9[42][4]}} & loc_sram_buff_w9[42][3:0]) | ({4{loc_sram_buff_w10[42][4]}} & loc_sram_buff_w10[42][3:0]) | ({4{loc_sram_buff_w11[42][4]}} & loc_sram_buff_w11[42][3:0]) | ({4{loc_sram_buff_w12[42][4]}} & loc_sram_buff_w12[42][3:0]) | ({4{loc_sram_buff_w13[42][4]}} & loc_sram_buff_w13[42][3:0]) | ({4{loc_sram_buff_w14[42][4]}} & loc_sram_buff_w14[42][3:0]) | ({4{loc_sram_buff_w15[42][4]}} & loc_sram_buff_w15[42][3:0]);
	loc_rdata_buff[ 851: 848] = ({4{loc_sram_buff_w0[43][4]}} & loc_sram_buff_w0[43][3:0]) | ({4{loc_sram_buff_w1[43][4]}} & loc_sram_buff_w1[43][3:0]) | ({4{loc_sram_buff_w2[43][4]}} & loc_sram_buff_w2[43][3:0]) | ({4{loc_sram_buff_w3[43][4]}} & loc_sram_buff_w3[43][3:0]) | ({4{loc_sram_buff_w4[43][4]}} & loc_sram_buff_w4[43][3:0]) | ({4{loc_sram_buff_w5[43][4]}} & loc_sram_buff_w5[43][3:0]) | ({4{loc_sram_buff_w6[43][4]}} & loc_sram_buff_w6[43][3:0]) | ({4{loc_sram_buff_w7[43][4]}} & loc_sram_buff_w7[43][3:0]) | ({4{loc_sram_buff_w8[43][4]}} & loc_sram_buff_w8[43][3:0]) | ({4{loc_sram_buff_w9[43][4]}} & loc_sram_buff_w9[43][3:0]) | ({4{loc_sram_buff_w10[43][4]}} & loc_sram_buff_w10[43][3:0]) | ({4{loc_sram_buff_w11[43][4]}} & loc_sram_buff_w11[43][3:0]) | ({4{loc_sram_buff_w12[43][4]}} & loc_sram_buff_w12[43][3:0]) | ({4{loc_sram_buff_w13[43][4]}} & loc_sram_buff_w13[43][3:0]) | ({4{loc_sram_buff_w14[43][4]}} & loc_sram_buff_w14[43][3:0]) | ({4{loc_sram_buff_w15[43][4]}} & loc_sram_buff_w15[43][3:0]);
	loc_rdata_buff[ 847: 844] = ({4{loc_sram_buff_w0[44][4]}} & loc_sram_buff_w0[44][3:0]) | ({4{loc_sram_buff_w1[44][4]}} & loc_sram_buff_w1[44][3:0]) | ({4{loc_sram_buff_w2[44][4]}} & loc_sram_buff_w2[44][3:0]) | ({4{loc_sram_buff_w3[44][4]}} & loc_sram_buff_w3[44][3:0]) | ({4{loc_sram_buff_w4[44][4]}} & loc_sram_buff_w4[44][3:0]) | ({4{loc_sram_buff_w5[44][4]}} & loc_sram_buff_w5[44][3:0]) | ({4{loc_sram_buff_w6[44][4]}} & loc_sram_buff_w6[44][3:0]) | ({4{loc_sram_buff_w7[44][4]}} & loc_sram_buff_w7[44][3:0]) | ({4{loc_sram_buff_w8[44][4]}} & loc_sram_buff_w8[44][3:0]) | ({4{loc_sram_buff_w9[44][4]}} & loc_sram_buff_w9[44][3:0]) | ({4{loc_sram_buff_w10[44][4]}} & loc_sram_buff_w10[44][3:0]) | ({4{loc_sram_buff_w11[44][4]}} & loc_sram_buff_w11[44][3:0]) | ({4{loc_sram_buff_w12[44][4]}} & loc_sram_buff_w12[44][3:0]) | ({4{loc_sram_buff_w13[44][4]}} & loc_sram_buff_w13[44][3:0]) | ({4{loc_sram_buff_w14[44][4]}} & loc_sram_buff_w14[44][3:0]) | ({4{loc_sram_buff_w15[44][4]}} & loc_sram_buff_w15[44][3:0]);
	loc_rdata_buff[ 843: 840] = ({4{loc_sram_buff_w0[45][4]}} & loc_sram_buff_w0[45][3:0]) | ({4{loc_sram_buff_w1[45][4]}} & loc_sram_buff_w1[45][3:0]) | ({4{loc_sram_buff_w2[45][4]}} & loc_sram_buff_w2[45][3:0]) | ({4{loc_sram_buff_w3[45][4]}} & loc_sram_buff_w3[45][3:0]) | ({4{loc_sram_buff_w4[45][4]}} & loc_sram_buff_w4[45][3:0]) | ({4{loc_sram_buff_w5[45][4]}} & loc_sram_buff_w5[45][3:0]) | ({4{loc_sram_buff_w6[45][4]}} & loc_sram_buff_w6[45][3:0]) | ({4{loc_sram_buff_w7[45][4]}} & loc_sram_buff_w7[45][3:0]) | ({4{loc_sram_buff_w8[45][4]}} & loc_sram_buff_w8[45][3:0]) | ({4{loc_sram_buff_w9[45][4]}} & loc_sram_buff_w9[45][3:0]) | ({4{loc_sram_buff_w10[45][4]}} & loc_sram_buff_w10[45][3:0]) | ({4{loc_sram_buff_w11[45][4]}} & loc_sram_buff_w11[45][3:0]) | ({4{loc_sram_buff_w12[45][4]}} & loc_sram_buff_w12[45][3:0]) | ({4{loc_sram_buff_w13[45][4]}} & loc_sram_buff_w13[45][3:0]) | ({4{loc_sram_buff_w14[45][4]}} & loc_sram_buff_w14[45][3:0]) | ({4{loc_sram_buff_w15[45][4]}} & loc_sram_buff_w15[45][3:0]);
	loc_rdata_buff[ 839: 836] = ({4{loc_sram_buff_w0[46][4]}} & loc_sram_buff_w0[46][3:0]) | ({4{loc_sram_buff_w1[46][4]}} & loc_sram_buff_w1[46][3:0]) | ({4{loc_sram_buff_w2[46][4]}} & loc_sram_buff_w2[46][3:0]) | ({4{loc_sram_buff_w3[46][4]}} & loc_sram_buff_w3[46][3:0]) | ({4{loc_sram_buff_w4[46][4]}} & loc_sram_buff_w4[46][3:0]) | ({4{loc_sram_buff_w5[46][4]}} & loc_sram_buff_w5[46][3:0]) | ({4{loc_sram_buff_w6[46][4]}} & loc_sram_buff_w6[46][3:0]) | ({4{loc_sram_buff_w7[46][4]}} & loc_sram_buff_w7[46][3:0]) | ({4{loc_sram_buff_w8[46][4]}} & loc_sram_buff_w8[46][3:0]) | ({4{loc_sram_buff_w9[46][4]}} & loc_sram_buff_w9[46][3:0]) | ({4{loc_sram_buff_w10[46][4]}} & loc_sram_buff_w10[46][3:0]) | ({4{loc_sram_buff_w11[46][4]}} & loc_sram_buff_w11[46][3:0]) | ({4{loc_sram_buff_w12[46][4]}} & loc_sram_buff_w12[46][3:0]) | ({4{loc_sram_buff_w13[46][4]}} & loc_sram_buff_w13[46][3:0]) | ({4{loc_sram_buff_w14[46][4]}} & loc_sram_buff_w14[46][3:0]) | ({4{loc_sram_buff_w15[46][4]}} & loc_sram_buff_w15[46][3:0]);
	loc_rdata_buff[ 835: 832] = ({4{loc_sram_buff_w0[47][4]}} & loc_sram_buff_w0[47][3:0]) | ({4{loc_sram_buff_w1[47][4]}} & loc_sram_buff_w1[47][3:0]) | ({4{loc_sram_buff_w2[47][4]}} & loc_sram_buff_w2[47][3:0]) | ({4{loc_sram_buff_w3[47][4]}} & loc_sram_buff_w3[47][3:0]) | ({4{loc_sram_buff_w4[47][4]}} & loc_sram_buff_w4[47][3:0]) | ({4{loc_sram_buff_w5[47][4]}} & loc_sram_buff_w5[47][3:0]) | ({4{loc_sram_buff_w6[47][4]}} & loc_sram_buff_w6[47][3:0]) | ({4{loc_sram_buff_w7[47][4]}} & loc_sram_buff_w7[47][3:0]) | ({4{loc_sram_buff_w8[47][4]}} & loc_sram_buff_w8[47][3:0]) | ({4{loc_sram_buff_w9[47][4]}} & loc_sram_buff_w9[47][3:0]) | ({4{loc_sram_buff_w10[47][4]}} & loc_sram_buff_w10[47][3:0]) | ({4{loc_sram_buff_w11[47][4]}} & loc_sram_buff_w11[47][3:0]) | ({4{loc_sram_buff_w12[47][4]}} & loc_sram_buff_w12[47][3:0]) | ({4{loc_sram_buff_w13[47][4]}} & loc_sram_buff_w13[47][3:0]) | ({4{loc_sram_buff_w14[47][4]}} & loc_sram_buff_w14[47][3:0]) | ({4{loc_sram_buff_w15[47][4]}} & loc_sram_buff_w15[47][3:0]);
	loc_rdata_buff[ 831: 828] = ({4{loc_sram_buff_w0[48][4]}} & loc_sram_buff_w0[48][3:0]) | ({4{loc_sram_buff_w1[48][4]}} & loc_sram_buff_w1[48][3:0]) | ({4{loc_sram_buff_w2[48][4]}} & loc_sram_buff_w2[48][3:0]) | ({4{loc_sram_buff_w3[48][4]}} & loc_sram_buff_w3[48][3:0]) | ({4{loc_sram_buff_w4[48][4]}} & loc_sram_buff_w4[48][3:0]) | ({4{loc_sram_buff_w5[48][4]}} & loc_sram_buff_w5[48][3:0]) | ({4{loc_sram_buff_w6[48][4]}} & loc_sram_buff_w6[48][3:0]) | ({4{loc_sram_buff_w7[48][4]}} & loc_sram_buff_w7[48][3:0]) | ({4{loc_sram_buff_w8[48][4]}} & loc_sram_buff_w8[48][3:0]) | ({4{loc_sram_buff_w9[48][4]}} & loc_sram_buff_w9[48][3:0]) | ({4{loc_sram_buff_w10[48][4]}} & loc_sram_buff_w10[48][3:0]) | ({4{loc_sram_buff_w11[48][4]}} & loc_sram_buff_w11[48][3:0]) | ({4{loc_sram_buff_w12[48][4]}} & loc_sram_buff_w12[48][3:0]) | ({4{loc_sram_buff_w13[48][4]}} & loc_sram_buff_w13[48][3:0]) | ({4{loc_sram_buff_w14[48][4]}} & loc_sram_buff_w14[48][3:0]) | ({4{loc_sram_buff_w15[48][4]}} & loc_sram_buff_w15[48][3:0]);
	loc_rdata_buff[ 827: 824] = ({4{loc_sram_buff_w0[49][4]}} & loc_sram_buff_w0[49][3:0]) | ({4{loc_sram_buff_w1[49][4]}} & loc_sram_buff_w1[49][3:0]) | ({4{loc_sram_buff_w2[49][4]}} & loc_sram_buff_w2[49][3:0]) | ({4{loc_sram_buff_w3[49][4]}} & loc_sram_buff_w3[49][3:0]) | ({4{loc_sram_buff_w4[49][4]}} & loc_sram_buff_w4[49][3:0]) | ({4{loc_sram_buff_w5[49][4]}} & loc_sram_buff_w5[49][3:0]) | ({4{loc_sram_buff_w6[49][4]}} & loc_sram_buff_w6[49][3:0]) | ({4{loc_sram_buff_w7[49][4]}} & loc_sram_buff_w7[49][3:0]) | ({4{loc_sram_buff_w8[49][4]}} & loc_sram_buff_w8[49][3:0]) | ({4{loc_sram_buff_w9[49][4]}} & loc_sram_buff_w9[49][3:0]) | ({4{loc_sram_buff_w10[49][4]}} & loc_sram_buff_w10[49][3:0]) | ({4{loc_sram_buff_w11[49][4]}} & loc_sram_buff_w11[49][3:0]) | ({4{loc_sram_buff_w12[49][4]}} & loc_sram_buff_w12[49][3:0]) | ({4{loc_sram_buff_w13[49][4]}} & loc_sram_buff_w13[49][3:0]) | ({4{loc_sram_buff_w14[49][4]}} & loc_sram_buff_w14[49][3:0]) | ({4{loc_sram_buff_w15[49][4]}} & loc_sram_buff_w15[49][3:0]);
	loc_rdata_buff[ 823: 820] = ({4{loc_sram_buff_w0[50][4]}} & loc_sram_buff_w0[50][3:0]) | ({4{loc_sram_buff_w1[50][4]}} & loc_sram_buff_w1[50][3:0]) | ({4{loc_sram_buff_w2[50][4]}} & loc_sram_buff_w2[50][3:0]) | ({4{loc_sram_buff_w3[50][4]}} & loc_sram_buff_w3[50][3:0]) | ({4{loc_sram_buff_w4[50][4]}} & loc_sram_buff_w4[50][3:0]) | ({4{loc_sram_buff_w5[50][4]}} & loc_sram_buff_w5[50][3:0]) | ({4{loc_sram_buff_w6[50][4]}} & loc_sram_buff_w6[50][3:0]) | ({4{loc_sram_buff_w7[50][4]}} & loc_sram_buff_w7[50][3:0]) | ({4{loc_sram_buff_w8[50][4]}} & loc_sram_buff_w8[50][3:0]) | ({4{loc_sram_buff_w9[50][4]}} & loc_sram_buff_w9[50][3:0]) | ({4{loc_sram_buff_w10[50][4]}} & loc_sram_buff_w10[50][3:0]) | ({4{loc_sram_buff_w11[50][4]}} & loc_sram_buff_w11[50][3:0]) | ({4{loc_sram_buff_w12[50][4]}} & loc_sram_buff_w12[50][3:0]) | ({4{loc_sram_buff_w13[50][4]}} & loc_sram_buff_w13[50][3:0]) | ({4{loc_sram_buff_w14[50][4]}} & loc_sram_buff_w14[50][3:0]) | ({4{loc_sram_buff_w15[50][4]}} & loc_sram_buff_w15[50][3:0]);
	loc_rdata_buff[ 819: 816] = ({4{loc_sram_buff_w0[51][4]}} & loc_sram_buff_w0[51][3:0]) | ({4{loc_sram_buff_w1[51][4]}} & loc_sram_buff_w1[51][3:0]) | ({4{loc_sram_buff_w2[51][4]}} & loc_sram_buff_w2[51][3:0]) | ({4{loc_sram_buff_w3[51][4]}} & loc_sram_buff_w3[51][3:0]) | ({4{loc_sram_buff_w4[51][4]}} & loc_sram_buff_w4[51][3:0]) | ({4{loc_sram_buff_w5[51][4]}} & loc_sram_buff_w5[51][3:0]) | ({4{loc_sram_buff_w6[51][4]}} & loc_sram_buff_w6[51][3:0]) | ({4{loc_sram_buff_w7[51][4]}} & loc_sram_buff_w7[51][3:0]) | ({4{loc_sram_buff_w8[51][4]}} & loc_sram_buff_w8[51][3:0]) | ({4{loc_sram_buff_w9[51][4]}} & loc_sram_buff_w9[51][3:0]) | ({4{loc_sram_buff_w10[51][4]}} & loc_sram_buff_w10[51][3:0]) | ({4{loc_sram_buff_w11[51][4]}} & loc_sram_buff_w11[51][3:0]) | ({4{loc_sram_buff_w12[51][4]}} & loc_sram_buff_w12[51][3:0]) | ({4{loc_sram_buff_w13[51][4]}} & loc_sram_buff_w13[51][3:0]) | ({4{loc_sram_buff_w14[51][4]}} & loc_sram_buff_w14[51][3:0]) | ({4{loc_sram_buff_w15[51][4]}} & loc_sram_buff_w15[51][3:0]);
	loc_rdata_buff[ 815: 812] = ({4{loc_sram_buff_w0[52][4]}} & loc_sram_buff_w0[52][3:0]) | ({4{loc_sram_buff_w1[52][4]}} & loc_sram_buff_w1[52][3:0]) | ({4{loc_sram_buff_w2[52][4]}} & loc_sram_buff_w2[52][3:0]) | ({4{loc_sram_buff_w3[52][4]}} & loc_sram_buff_w3[52][3:0]) | ({4{loc_sram_buff_w4[52][4]}} & loc_sram_buff_w4[52][3:0]) | ({4{loc_sram_buff_w5[52][4]}} & loc_sram_buff_w5[52][3:0]) | ({4{loc_sram_buff_w6[52][4]}} & loc_sram_buff_w6[52][3:0]) | ({4{loc_sram_buff_w7[52][4]}} & loc_sram_buff_w7[52][3:0]) | ({4{loc_sram_buff_w8[52][4]}} & loc_sram_buff_w8[52][3:0]) | ({4{loc_sram_buff_w9[52][4]}} & loc_sram_buff_w9[52][3:0]) | ({4{loc_sram_buff_w10[52][4]}} & loc_sram_buff_w10[52][3:0]) | ({4{loc_sram_buff_w11[52][4]}} & loc_sram_buff_w11[52][3:0]) | ({4{loc_sram_buff_w12[52][4]}} & loc_sram_buff_w12[52][3:0]) | ({4{loc_sram_buff_w13[52][4]}} & loc_sram_buff_w13[52][3:0]) | ({4{loc_sram_buff_w14[52][4]}} & loc_sram_buff_w14[52][3:0]) | ({4{loc_sram_buff_w15[52][4]}} & loc_sram_buff_w15[52][3:0]);
	loc_rdata_buff[ 811: 808] = ({4{loc_sram_buff_w0[53][4]}} & loc_sram_buff_w0[53][3:0]) | ({4{loc_sram_buff_w1[53][4]}} & loc_sram_buff_w1[53][3:0]) | ({4{loc_sram_buff_w2[53][4]}} & loc_sram_buff_w2[53][3:0]) | ({4{loc_sram_buff_w3[53][4]}} & loc_sram_buff_w3[53][3:0]) | ({4{loc_sram_buff_w4[53][4]}} & loc_sram_buff_w4[53][3:0]) | ({4{loc_sram_buff_w5[53][4]}} & loc_sram_buff_w5[53][3:0]) | ({4{loc_sram_buff_w6[53][4]}} & loc_sram_buff_w6[53][3:0]) | ({4{loc_sram_buff_w7[53][4]}} & loc_sram_buff_w7[53][3:0]) | ({4{loc_sram_buff_w8[53][4]}} & loc_sram_buff_w8[53][3:0]) | ({4{loc_sram_buff_w9[53][4]}} & loc_sram_buff_w9[53][3:0]) | ({4{loc_sram_buff_w10[53][4]}} & loc_sram_buff_w10[53][3:0]) | ({4{loc_sram_buff_w11[53][4]}} & loc_sram_buff_w11[53][3:0]) | ({4{loc_sram_buff_w12[53][4]}} & loc_sram_buff_w12[53][3:0]) | ({4{loc_sram_buff_w13[53][4]}} & loc_sram_buff_w13[53][3:0]) | ({4{loc_sram_buff_w14[53][4]}} & loc_sram_buff_w14[53][3:0]) | ({4{loc_sram_buff_w15[53][4]}} & loc_sram_buff_w15[53][3:0]);
	loc_rdata_buff[ 807: 804] = ({4{loc_sram_buff_w0[54][4]}} & loc_sram_buff_w0[54][3:0]) | ({4{loc_sram_buff_w1[54][4]}} & loc_sram_buff_w1[54][3:0]) | ({4{loc_sram_buff_w2[54][4]}} & loc_sram_buff_w2[54][3:0]) | ({4{loc_sram_buff_w3[54][4]}} & loc_sram_buff_w3[54][3:0]) | ({4{loc_sram_buff_w4[54][4]}} & loc_sram_buff_w4[54][3:0]) | ({4{loc_sram_buff_w5[54][4]}} & loc_sram_buff_w5[54][3:0]) | ({4{loc_sram_buff_w6[54][4]}} & loc_sram_buff_w6[54][3:0]) | ({4{loc_sram_buff_w7[54][4]}} & loc_sram_buff_w7[54][3:0]) | ({4{loc_sram_buff_w8[54][4]}} & loc_sram_buff_w8[54][3:0]) | ({4{loc_sram_buff_w9[54][4]}} & loc_sram_buff_w9[54][3:0]) | ({4{loc_sram_buff_w10[54][4]}} & loc_sram_buff_w10[54][3:0]) | ({4{loc_sram_buff_w11[54][4]}} & loc_sram_buff_w11[54][3:0]) | ({4{loc_sram_buff_w12[54][4]}} & loc_sram_buff_w12[54][3:0]) | ({4{loc_sram_buff_w13[54][4]}} & loc_sram_buff_w13[54][3:0]) | ({4{loc_sram_buff_w14[54][4]}} & loc_sram_buff_w14[54][3:0]) | ({4{loc_sram_buff_w15[54][4]}} & loc_sram_buff_w15[54][3:0]);
	loc_rdata_buff[ 803: 800] = ({4{loc_sram_buff_w0[55][4]}} & loc_sram_buff_w0[55][3:0]) | ({4{loc_sram_buff_w1[55][4]}} & loc_sram_buff_w1[55][3:0]) | ({4{loc_sram_buff_w2[55][4]}} & loc_sram_buff_w2[55][3:0]) | ({4{loc_sram_buff_w3[55][4]}} & loc_sram_buff_w3[55][3:0]) | ({4{loc_sram_buff_w4[55][4]}} & loc_sram_buff_w4[55][3:0]) | ({4{loc_sram_buff_w5[55][4]}} & loc_sram_buff_w5[55][3:0]) | ({4{loc_sram_buff_w6[55][4]}} & loc_sram_buff_w6[55][3:0]) | ({4{loc_sram_buff_w7[55][4]}} & loc_sram_buff_w7[55][3:0]) | ({4{loc_sram_buff_w8[55][4]}} & loc_sram_buff_w8[55][3:0]) | ({4{loc_sram_buff_w9[55][4]}} & loc_sram_buff_w9[55][3:0]) | ({4{loc_sram_buff_w10[55][4]}} & loc_sram_buff_w10[55][3:0]) | ({4{loc_sram_buff_w11[55][4]}} & loc_sram_buff_w11[55][3:0]) | ({4{loc_sram_buff_w12[55][4]}} & loc_sram_buff_w12[55][3:0]) | ({4{loc_sram_buff_w13[55][4]}} & loc_sram_buff_w13[55][3:0]) | ({4{loc_sram_buff_w14[55][4]}} & loc_sram_buff_w14[55][3:0]) | ({4{loc_sram_buff_w15[55][4]}} & loc_sram_buff_w15[55][3:0]);
	loc_rdata_buff[ 799: 796] = ({4{loc_sram_buff_w0[56][4]}} & loc_sram_buff_w0[56][3:0]) | ({4{loc_sram_buff_w1[56][4]}} & loc_sram_buff_w1[56][3:0]) | ({4{loc_sram_buff_w2[56][4]}} & loc_sram_buff_w2[56][3:0]) | ({4{loc_sram_buff_w3[56][4]}} & loc_sram_buff_w3[56][3:0]) | ({4{loc_sram_buff_w4[56][4]}} & loc_sram_buff_w4[56][3:0]) | ({4{loc_sram_buff_w5[56][4]}} & loc_sram_buff_w5[56][3:0]) | ({4{loc_sram_buff_w6[56][4]}} & loc_sram_buff_w6[56][3:0]) | ({4{loc_sram_buff_w7[56][4]}} & loc_sram_buff_w7[56][3:0]) | ({4{loc_sram_buff_w8[56][4]}} & loc_sram_buff_w8[56][3:0]) | ({4{loc_sram_buff_w9[56][4]}} & loc_sram_buff_w9[56][3:0]) | ({4{loc_sram_buff_w10[56][4]}} & loc_sram_buff_w10[56][3:0]) | ({4{loc_sram_buff_w11[56][4]}} & loc_sram_buff_w11[56][3:0]) | ({4{loc_sram_buff_w12[56][4]}} & loc_sram_buff_w12[56][3:0]) | ({4{loc_sram_buff_w13[56][4]}} & loc_sram_buff_w13[56][3:0]) | ({4{loc_sram_buff_w14[56][4]}} & loc_sram_buff_w14[56][3:0]) | ({4{loc_sram_buff_w15[56][4]}} & loc_sram_buff_w15[56][3:0]);
	loc_rdata_buff[ 795: 792] = ({4{loc_sram_buff_w0[57][4]}} & loc_sram_buff_w0[57][3:0]) | ({4{loc_sram_buff_w1[57][4]}} & loc_sram_buff_w1[57][3:0]) | ({4{loc_sram_buff_w2[57][4]}} & loc_sram_buff_w2[57][3:0]) | ({4{loc_sram_buff_w3[57][4]}} & loc_sram_buff_w3[57][3:0]) | ({4{loc_sram_buff_w4[57][4]}} & loc_sram_buff_w4[57][3:0]) | ({4{loc_sram_buff_w5[57][4]}} & loc_sram_buff_w5[57][3:0]) | ({4{loc_sram_buff_w6[57][4]}} & loc_sram_buff_w6[57][3:0]) | ({4{loc_sram_buff_w7[57][4]}} & loc_sram_buff_w7[57][3:0]) | ({4{loc_sram_buff_w8[57][4]}} & loc_sram_buff_w8[57][3:0]) | ({4{loc_sram_buff_w9[57][4]}} & loc_sram_buff_w9[57][3:0]) | ({4{loc_sram_buff_w10[57][4]}} & loc_sram_buff_w10[57][3:0]) | ({4{loc_sram_buff_w11[57][4]}} & loc_sram_buff_w11[57][3:0]) | ({4{loc_sram_buff_w12[57][4]}} & loc_sram_buff_w12[57][3:0]) | ({4{loc_sram_buff_w13[57][4]}} & loc_sram_buff_w13[57][3:0]) | ({4{loc_sram_buff_w14[57][4]}} & loc_sram_buff_w14[57][3:0]) | ({4{loc_sram_buff_w15[57][4]}} & loc_sram_buff_w15[57][3:0]);
	loc_rdata_buff[ 791: 788] = ({4{loc_sram_buff_w0[58][4]}} & loc_sram_buff_w0[58][3:0]) | ({4{loc_sram_buff_w1[58][4]}} & loc_sram_buff_w1[58][3:0]) | ({4{loc_sram_buff_w2[58][4]}} & loc_sram_buff_w2[58][3:0]) | ({4{loc_sram_buff_w3[58][4]}} & loc_sram_buff_w3[58][3:0]) | ({4{loc_sram_buff_w4[58][4]}} & loc_sram_buff_w4[58][3:0]) | ({4{loc_sram_buff_w5[58][4]}} & loc_sram_buff_w5[58][3:0]) | ({4{loc_sram_buff_w6[58][4]}} & loc_sram_buff_w6[58][3:0]) | ({4{loc_sram_buff_w7[58][4]}} & loc_sram_buff_w7[58][3:0]) | ({4{loc_sram_buff_w8[58][4]}} & loc_sram_buff_w8[58][3:0]) | ({4{loc_sram_buff_w9[58][4]}} & loc_sram_buff_w9[58][3:0]) | ({4{loc_sram_buff_w10[58][4]}} & loc_sram_buff_w10[58][3:0]) | ({4{loc_sram_buff_w11[58][4]}} & loc_sram_buff_w11[58][3:0]) | ({4{loc_sram_buff_w12[58][4]}} & loc_sram_buff_w12[58][3:0]) | ({4{loc_sram_buff_w13[58][4]}} & loc_sram_buff_w13[58][3:0]) | ({4{loc_sram_buff_w14[58][4]}} & loc_sram_buff_w14[58][3:0]) | ({4{loc_sram_buff_w15[58][4]}} & loc_sram_buff_w15[58][3:0]);
	loc_rdata_buff[ 787: 784] = ({4{loc_sram_buff_w0[59][4]}} & loc_sram_buff_w0[59][3:0]) | ({4{loc_sram_buff_w1[59][4]}} & loc_sram_buff_w1[59][3:0]) | ({4{loc_sram_buff_w2[59][4]}} & loc_sram_buff_w2[59][3:0]) | ({4{loc_sram_buff_w3[59][4]}} & loc_sram_buff_w3[59][3:0]) | ({4{loc_sram_buff_w4[59][4]}} & loc_sram_buff_w4[59][3:0]) | ({4{loc_sram_buff_w5[59][4]}} & loc_sram_buff_w5[59][3:0]) | ({4{loc_sram_buff_w6[59][4]}} & loc_sram_buff_w6[59][3:0]) | ({4{loc_sram_buff_w7[59][4]}} & loc_sram_buff_w7[59][3:0]) | ({4{loc_sram_buff_w8[59][4]}} & loc_sram_buff_w8[59][3:0]) | ({4{loc_sram_buff_w9[59][4]}} & loc_sram_buff_w9[59][3:0]) | ({4{loc_sram_buff_w10[59][4]}} & loc_sram_buff_w10[59][3:0]) | ({4{loc_sram_buff_w11[59][4]}} & loc_sram_buff_w11[59][3:0]) | ({4{loc_sram_buff_w12[59][4]}} & loc_sram_buff_w12[59][3:0]) | ({4{loc_sram_buff_w13[59][4]}} & loc_sram_buff_w13[59][3:0]) | ({4{loc_sram_buff_w14[59][4]}} & loc_sram_buff_w14[59][3:0]) | ({4{loc_sram_buff_w15[59][4]}} & loc_sram_buff_w15[59][3:0]);
	loc_rdata_buff[ 783: 780] = ({4{loc_sram_buff_w0[60][4]}} & loc_sram_buff_w0[60][3:0]) | ({4{loc_sram_buff_w1[60][4]}} & loc_sram_buff_w1[60][3:0]) | ({4{loc_sram_buff_w2[60][4]}} & loc_sram_buff_w2[60][3:0]) | ({4{loc_sram_buff_w3[60][4]}} & loc_sram_buff_w3[60][3:0]) | ({4{loc_sram_buff_w4[60][4]}} & loc_sram_buff_w4[60][3:0]) | ({4{loc_sram_buff_w5[60][4]}} & loc_sram_buff_w5[60][3:0]) | ({4{loc_sram_buff_w6[60][4]}} & loc_sram_buff_w6[60][3:0]) | ({4{loc_sram_buff_w7[60][4]}} & loc_sram_buff_w7[60][3:0]) | ({4{loc_sram_buff_w8[60][4]}} & loc_sram_buff_w8[60][3:0]) | ({4{loc_sram_buff_w9[60][4]}} & loc_sram_buff_w9[60][3:0]) | ({4{loc_sram_buff_w10[60][4]}} & loc_sram_buff_w10[60][3:0]) | ({4{loc_sram_buff_w11[60][4]}} & loc_sram_buff_w11[60][3:0]) | ({4{loc_sram_buff_w12[60][4]}} & loc_sram_buff_w12[60][3:0]) | ({4{loc_sram_buff_w13[60][4]}} & loc_sram_buff_w13[60][3:0]) | ({4{loc_sram_buff_w14[60][4]}} & loc_sram_buff_w14[60][3:0]) | ({4{loc_sram_buff_w15[60][4]}} & loc_sram_buff_w15[60][3:0]);
	loc_rdata_buff[ 779: 776] = ({4{loc_sram_buff_w0[61][4]}} & loc_sram_buff_w0[61][3:0]) | ({4{loc_sram_buff_w1[61][4]}} & loc_sram_buff_w1[61][3:0]) | ({4{loc_sram_buff_w2[61][4]}} & loc_sram_buff_w2[61][3:0]) | ({4{loc_sram_buff_w3[61][4]}} & loc_sram_buff_w3[61][3:0]) | ({4{loc_sram_buff_w4[61][4]}} & loc_sram_buff_w4[61][3:0]) | ({4{loc_sram_buff_w5[61][4]}} & loc_sram_buff_w5[61][3:0]) | ({4{loc_sram_buff_w6[61][4]}} & loc_sram_buff_w6[61][3:0]) | ({4{loc_sram_buff_w7[61][4]}} & loc_sram_buff_w7[61][3:0]) | ({4{loc_sram_buff_w8[61][4]}} & loc_sram_buff_w8[61][3:0]) | ({4{loc_sram_buff_w9[61][4]}} & loc_sram_buff_w9[61][3:0]) | ({4{loc_sram_buff_w10[61][4]}} & loc_sram_buff_w10[61][3:0]) | ({4{loc_sram_buff_w11[61][4]}} & loc_sram_buff_w11[61][3:0]) | ({4{loc_sram_buff_w12[61][4]}} & loc_sram_buff_w12[61][3:0]) | ({4{loc_sram_buff_w13[61][4]}} & loc_sram_buff_w13[61][3:0]) | ({4{loc_sram_buff_w14[61][4]}} & loc_sram_buff_w14[61][3:0]) | ({4{loc_sram_buff_w15[61][4]}} & loc_sram_buff_w15[61][3:0]);
	loc_rdata_buff[ 775: 772] = ({4{loc_sram_buff_w0[62][4]}} & loc_sram_buff_w0[62][3:0]) | ({4{loc_sram_buff_w1[62][4]}} & loc_sram_buff_w1[62][3:0]) | ({4{loc_sram_buff_w2[62][4]}} & loc_sram_buff_w2[62][3:0]) | ({4{loc_sram_buff_w3[62][4]}} & loc_sram_buff_w3[62][3:0]) | ({4{loc_sram_buff_w4[62][4]}} & loc_sram_buff_w4[62][3:0]) | ({4{loc_sram_buff_w5[62][4]}} & loc_sram_buff_w5[62][3:0]) | ({4{loc_sram_buff_w6[62][4]}} & loc_sram_buff_w6[62][3:0]) | ({4{loc_sram_buff_w7[62][4]}} & loc_sram_buff_w7[62][3:0]) | ({4{loc_sram_buff_w8[62][4]}} & loc_sram_buff_w8[62][3:0]) | ({4{loc_sram_buff_w9[62][4]}} & loc_sram_buff_w9[62][3:0]) | ({4{loc_sram_buff_w10[62][4]}} & loc_sram_buff_w10[62][3:0]) | ({4{loc_sram_buff_w11[62][4]}} & loc_sram_buff_w11[62][3:0]) | ({4{loc_sram_buff_w12[62][4]}} & loc_sram_buff_w12[62][3:0]) | ({4{loc_sram_buff_w13[62][4]}} & loc_sram_buff_w13[62][3:0]) | ({4{loc_sram_buff_w14[62][4]}} & loc_sram_buff_w14[62][3:0]) | ({4{loc_sram_buff_w15[62][4]}} & loc_sram_buff_w15[62][3:0]);
	loc_rdata_buff[ 771: 768] = ({4{loc_sram_buff_w0[63][4]}} & loc_sram_buff_w0[63][3:0]) | ({4{loc_sram_buff_w1[63][4]}} & loc_sram_buff_w1[63][3:0]) | ({4{loc_sram_buff_w2[63][4]}} & loc_sram_buff_w2[63][3:0]) | ({4{loc_sram_buff_w3[63][4]}} & loc_sram_buff_w3[63][3:0]) | ({4{loc_sram_buff_w4[63][4]}} & loc_sram_buff_w4[63][3:0]) | ({4{loc_sram_buff_w5[63][4]}} & loc_sram_buff_w5[63][3:0]) | ({4{loc_sram_buff_w6[63][4]}} & loc_sram_buff_w6[63][3:0]) | ({4{loc_sram_buff_w7[63][4]}} & loc_sram_buff_w7[63][3:0]) | ({4{loc_sram_buff_w8[63][4]}} & loc_sram_buff_w8[63][3:0]) | ({4{loc_sram_buff_w9[63][4]}} & loc_sram_buff_w9[63][3:0]) | ({4{loc_sram_buff_w10[63][4]}} & loc_sram_buff_w10[63][3:0]) | ({4{loc_sram_buff_w11[63][4]}} & loc_sram_buff_w11[63][3:0]) | ({4{loc_sram_buff_w12[63][4]}} & loc_sram_buff_w12[63][3:0]) | ({4{loc_sram_buff_w13[63][4]}} & loc_sram_buff_w13[63][3:0]) | ({4{loc_sram_buff_w14[63][4]}} & loc_sram_buff_w14[63][3:0]) | ({4{loc_sram_buff_w15[63][4]}} & loc_sram_buff_w15[63][3:0]);
	loc_rdata_buff[ 767: 764] = ({4{loc_sram_buff_w0[64][4]}} & loc_sram_buff_w0[64][3:0]) | ({4{loc_sram_buff_w1[64][4]}} & loc_sram_buff_w1[64][3:0]) | ({4{loc_sram_buff_w2[64][4]}} & loc_sram_buff_w2[64][3:0]) | ({4{loc_sram_buff_w3[64][4]}} & loc_sram_buff_w3[64][3:0]) | ({4{loc_sram_buff_w4[64][4]}} & loc_sram_buff_w4[64][3:0]) | ({4{loc_sram_buff_w5[64][4]}} & loc_sram_buff_w5[64][3:0]) | ({4{loc_sram_buff_w6[64][4]}} & loc_sram_buff_w6[64][3:0]) | ({4{loc_sram_buff_w7[64][4]}} & loc_sram_buff_w7[64][3:0]) | ({4{loc_sram_buff_w8[64][4]}} & loc_sram_buff_w8[64][3:0]) | ({4{loc_sram_buff_w9[64][4]}} & loc_sram_buff_w9[64][3:0]) | ({4{loc_sram_buff_w10[64][4]}} & loc_sram_buff_w10[64][3:0]) | ({4{loc_sram_buff_w11[64][4]}} & loc_sram_buff_w11[64][3:0]) | ({4{loc_sram_buff_w12[64][4]}} & loc_sram_buff_w12[64][3:0]) | ({4{loc_sram_buff_w13[64][4]}} & loc_sram_buff_w13[64][3:0]) | ({4{loc_sram_buff_w14[64][4]}} & loc_sram_buff_w14[64][3:0]) | ({4{loc_sram_buff_w15[64][4]}} & loc_sram_buff_w15[64][3:0]);
	loc_rdata_buff[ 763: 760] = ({4{loc_sram_buff_w0[65][4]}} & loc_sram_buff_w0[65][3:0]) | ({4{loc_sram_buff_w1[65][4]}} & loc_sram_buff_w1[65][3:0]) | ({4{loc_sram_buff_w2[65][4]}} & loc_sram_buff_w2[65][3:0]) | ({4{loc_sram_buff_w3[65][4]}} & loc_sram_buff_w3[65][3:0]) | ({4{loc_sram_buff_w4[65][4]}} & loc_sram_buff_w4[65][3:0]) | ({4{loc_sram_buff_w5[65][4]}} & loc_sram_buff_w5[65][3:0]) | ({4{loc_sram_buff_w6[65][4]}} & loc_sram_buff_w6[65][3:0]) | ({4{loc_sram_buff_w7[65][4]}} & loc_sram_buff_w7[65][3:0]) | ({4{loc_sram_buff_w8[65][4]}} & loc_sram_buff_w8[65][3:0]) | ({4{loc_sram_buff_w9[65][4]}} & loc_sram_buff_w9[65][3:0]) | ({4{loc_sram_buff_w10[65][4]}} & loc_sram_buff_w10[65][3:0]) | ({4{loc_sram_buff_w11[65][4]}} & loc_sram_buff_w11[65][3:0]) | ({4{loc_sram_buff_w12[65][4]}} & loc_sram_buff_w12[65][3:0]) | ({4{loc_sram_buff_w13[65][4]}} & loc_sram_buff_w13[65][3:0]) | ({4{loc_sram_buff_w14[65][4]}} & loc_sram_buff_w14[65][3:0]) | ({4{loc_sram_buff_w15[65][4]}} & loc_sram_buff_w15[65][3:0]);
	loc_rdata_buff[ 759: 756] = ({4{loc_sram_buff_w0[66][4]}} & loc_sram_buff_w0[66][3:0]) | ({4{loc_sram_buff_w1[66][4]}} & loc_sram_buff_w1[66][3:0]) | ({4{loc_sram_buff_w2[66][4]}} & loc_sram_buff_w2[66][3:0]) | ({4{loc_sram_buff_w3[66][4]}} & loc_sram_buff_w3[66][3:0]) | ({4{loc_sram_buff_w4[66][4]}} & loc_sram_buff_w4[66][3:0]) | ({4{loc_sram_buff_w5[66][4]}} & loc_sram_buff_w5[66][3:0]) | ({4{loc_sram_buff_w6[66][4]}} & loc_sram_buff_w6[66][3:0]) | ({4{loc_sram_buff_w7[66][4]}} & loc_sram_buff_w7[66][3:0]) | ({4{loc_sram_buff_w8[66][4]}} & loc_sram_buff_w8[66][3:0]) | ({4{loc_sram_buff_w9[66][4]}} & loc_sram_buff_w9[66][3:0]) | ({4{loc_sram_buff_w10[66][4]}} & loc_sram_buff_w10[66][3:0]) | ({4{loc_sram_buff_w11[66][4]}} & loc_sram_buff_w11[66][3:0]) | ({4{loc_sram_buff_w12[66][4]}} & loc_sram_buff_w12[66][3:0]) | ({4{loc_sram_buff_w13[66][4]}} & loc_sram_buff_w13[66][3:0]) | ({4{loc_sram_buff_w14[66][4]}} & loc_sram_buff_w14[66][3:0]) | ({4{loc_sram_buff_w15[66][4]}} & loc_sram_buff_w15[66][3:0]);
	loc_rdata_buff[ 755: 752] = ({4{loc_sram_buff_w0[67][4]}} & loc_sram_buff_w0[67][3:0]) | ({4{loc_sram_buff_w1[67][4]}} & loc_sram_buff_w1[67][3:0]) | ({4{loc_sram_buff_w2[67][4]}} & loc_sram_buff_w2[67][3:0]) | ({4{loc_sram_buff_w3[67][4]}} & loc_sram_buff_w3[67][3:0]) | ({4{loc_sram_buff_w4[67][4]}} & loc_sram_buff_w4[67][3:0]) | ({4{loc_sram_buff_w5[67][4]}} & loc_sram_buff_w5[67][3:0]) | ({4{loc_sram_buff_w6[67][4]}} & loc_sram_buff_w6[67][3:0]) | ({4{loc_sram_buff_w7[67][4]}} & loc_sram_buff_w7[67][3:0]) | ({4{loc_sram_buff_w8[67][4]}} & loc_sram_buff_w8[67][3:0]) | ({4{loc_sram_buff_w9[67][4]}} & loc_sram_buff_w9[67][3:0]) | ({4{loc_sram_buff_w10[67][4]}} & loc_sram_buff_w10[67][3:0]) | ({4{loc_sram_buff_w11[67][4]}} & loc_sram_buff_w11[67][3:0]) | ({4{loc_sram_buff_w12[67][4]}} & loc_sram_buff_w12[67][3:0]) | ({4{loc_sram_buff_w13[67][4]}} & loc_sram_buff_w13[67][3:0]) | ({4{loc_sram_buff_w14[67][4]}} & loc_sram_buff_w14[67][3:0]) | ({4{loc_sram_buff_w15[67][4]}} & loc_sram_buff_w15[67][3:0]);
	loc_rdata_buff[ 751: 748] = ({4{loc_sram_buff_w0[68][4]}} & loc_sram_buff_w0[68][3:0]) | ({4{loc_sram_buff_w1[68][4]}} & loc_sram_buff_w1[68][3:0]) | ({4{loc_sram_buff_w2[68][4]}} & loc_sram_buff_w2[68][3:0]) | ({4{loc_sram_buff_w3[68][4]}} & loc_sram_buff_w3[68][3:0]) | ({4{loc_sram_buff_w4[68][4]}} & loc_sram_buff_w4[68][3:0]) | ({4{loc_sram_buff_w5[68][4]}} & loc_sram_buff_w5[68][3:0]) | ({4{loc_sram_buff_w6[68][4]}} & loc_sram_buff_w6[68][3:0]) | ({4{loc_sram_buff_w7[68][4]}} & loc_sram_buff_w7[68][3:0]) | ({4{loc_sram_buff_w8[68][4]}} & loc_sram_buff_w8[68][3:0]) | ({4{loc_sram_buff_w9[68][4]}} & loc_sram_buff_w9[68][3:0]) | ({4{loc_sram_buff_w10[68][4]}} & loc_sram_buff_w10[68][3:0]) | ({4{loc_sram_buff_w11[68][4]}} & loc_sram_buff_w11[68][3:0]) | ({4{loc_sram_buff_w12[68][4]}} & loc_sram_buff_w12[68][3:0]) | ({4{loc_sram_buff_w13[68][4]}} & loc_sram_buff_w13[68][3:0]) | ({4{loc_sram_buff_w14[68][4]}} & loc_sram_buff_w14[68][3:0]) | ({4{loc_sram_buff_w15[68][4]}} & loc_sram_buff_w15[68][3:0]);
	loc_rdata_buff[ 747: 744] = ({4{loc_sram_buff_w0[69][4]}} & loc_sram_buff_w0[69][3:0]) | ({4{loc_sram_buff_w1[69][4]}} & loc_sram_buff_w1[69][3:0]) | ({4{loc_sram_buff_w2[69][4]}} & loc_sram_buff_w2[69][3:0]) | ({4{loc_sram_buff_w3[69][4]}} & loc_sram_buff_w3[69][3:0]) | ({4{loc_sram_buff_w4[69][4]}} & loc_sram_buff_w4[69][3:0]) | ({4{loc_sram_buff_w5[69][4]}} & loc_sram_buff_w5[69][3:0]) | ({4{loc_sram_buff_w6[69][4]}} & loc_sram_buff_w6[69][3:0]) | ({4{loc_sram_buff_w7[69][4]}} & loc_sram_buff_w7[69][3:0]) | ({4{loc_sram_buff_w8[69][4]}} & loc_sram_buff_w8[69][3:0]) | ({4{loc_sram_buff_w9[69][4]}} & loc_sram_buff_w9[69][3:0]) | ({4{loc_sram_buff_w10[69][4]}} & loc_sram_buff_w10[69][3:0]) | ({4{loc_sram_buff_w11[69][4]}} & loc_sram_buff_w11[69][3:0]) | ({4{loc_sram_buff_w12[69][4]}} & loc_sram_buff_w12[69][3:0]) | ({4{loc_sram_buff_w13[69][4]}} & loc_sram_buff_w13[69][3:0]) | ({4{loc_sram_buff_w14[69][4]}} & loc_sram_buff_w14[69][3:0]) | ({4{loc_sram_buff_w15[69][4]}} & loc_sram_buff_w15[69][3:0]);
	loc_rdata_buff[ 743: 740] = ({4{loc_sram_buff_w0[70][4]}} & loc_sram_buff_w0[70][3:0]) | ({4{loc_sram_buff_w1[70][4]}} & loc_sram_buff_w1[70][3:0]) | ({4{loc_sram_buff_w2[70][4]}} & loc_sram_buff_w2[70][3:0]) | ({4{loc_sram_buff_w3[70][4]}} & loc_sram_buff_w3[70][3:0]) | ({4{loc_sram_buff_w4[70][4]}} & loc_sram_buff_w4[70][3:0]) | ({4{loc_sram_buff_w5[70][4]}} & loc_sram_buff_w5[70][3:0]) | ({4{loc_sram_buff_w6[70][4]}} & loc_sram_buff_w6[70][3:0]) | ({4{loc_sram_buff_w7[70][4]}} & loc_sram_buff_w7[70][3:0]) | ({4{loc_sram_buff_w8[70][4]}} & loc_sram_buff_w8[70][3:0]) | ({4{loc_sram_buff_w9[70][4]}} & loc_sram_buff_w9[70][3:0]) | ({4{loc_sram_buff_w10[70][4]}} & loc_sram_buff_w10[70][3:0]) | ({4{loc_sram_buff_w11[70][4]}} & loc_sram_buff_w11[70][3:0]) | ({4{loc_sram_buff_w12[70][4]}} & loc_sram_buff_w12[70][3:0]) | ({4{loc_sram_buff_w13[70][4]}} & loc_sram_buff_w13[70][3:0]) | ({4{loc_sram_buff_w14[70][4]}} & loc_sram_buff_w14[70][3:0]) | ({4{loc_sram_buff_w15[70][4]}} & loc_sram_buff_w15[70][3:0]);
	loc_rdata_buff[ 739: 736] = ({4{loc_sram_buff_w0[71][4]}} & loc_sram_buff_w0[71][3:0]) | ({4{loc_sram_buff_w1[71][4]}} & loc_sram_buff_w1[71][3:0]) | ({4{loc_sram_buff_w2[71][4]}} & loc_sram_buff_w2[71][3:0]) | ({4{loc_sram_buff_w3[71][4]}} & loc_sram_buff_w3[71][3:0]) | ({4{loc_sram_buff_w4[71][4]}} & loc_sram_buff_w4[71][3:0]) | ({4{loc_sram_buff_w5[71][4]}} & loc_sram_buff_w5[71][3:0]) | ({4{loc_sram_buff_w6[71][4]}} & loc_sram_buff_w6[71][3:0]) | ({4{loc_sram_buff_w7[71][4]}} & loc_sram_buff_w7[71][3:0]) | ({4{loc_sram_buff_w8[71][4]}} & loc_sram_buff_w8[71][3:0]) | ({4{loc_sram_buff_w9[71][4]}} & loc_sram_buff_w9[71][3:0]) | ({4{loc_sram_buff_w10[71][4]}} & loc_sram_buff_w10[71][3:0]) | ({4{loc_sram_buff_w11[71][4]}} & loc_sram_buff_w11[71][3:0]) | ({4{loc_sram_buff_w12[71][4]}} & loc_sram_buff_w12[71][3:0]) | ({4{loc_sram_buff_w13[71][4]}} & loc_sram_buff_w13[71][3:0]) | ({4{loc_sram_buff_w14[71][4]}} & loc_sram_buff_w14[71][3:0]) | ({4{loc_sram_buff_w15[71][4]}} & loc_sram_buff_w15[71][3:0]);
	loc_rdata_buff[ 735: 732] = ({4{loc_sram_buff_w0[72][4]}} & loc_sram_buff_w0[72][3:0]) | ({4{loc_sram_buff_w1[72][4]}} & loc_sram_buff_w1[72][3:0]) | ({4{loc_sram_buff_w2[72][4]}} & loc_sram_buff_w2[72][3:0]) | ({4{loc_sram_buff_w3[72][4]}} & loc_sram_buff_w3[72][3:0]) | ({4{loc_sram_buff_w4[72][4]}} & loc_sram_buff_w4[72][3:0]) | ({4{loc_sram_buff_w5[72][4]}} & loc_sram_buff_w5[72][3:0]) | ({4{loc_sram_buff_w6[72][4]}} & loc_sram_buff_w6[72][3:0]) | ({4{loc_sram_buff_w7[72][4]}} & loc_sram_buff_w7[72][3:0]) | ({4{loc_sram_buff_w8[72][4]}} & loc_sram_buff_w8[72][3:0]) | ({4{loc_sram_buff_w9[72][4]}} & loc_sram_buff_w9[72][3:0]) | ({4{loc_sram_buff_w10[72][4]}} & loc_sram_buff_w10[72][3:0]) | ({4{loc_sram_buff_w11[72][4]}} & loc_sram_buff_w11[72][3:0]) | ({4{loc_sram_buff_w12[72][4]}} & loc_sram_buff_w12[72][3:0]) | ({4{loc_sram_buff_w13[72][4]}} & loc_sram_buff_w13[72][3:0]) | ({4{loc_sram_buff_w14[72][4]}} & loc_sram_buff_w14[72][3:0]) | ({4{loc_sram_buff_w15[72][4]}} & loc_sram_buff_w15[72][3:0]);
	loc_rdata_buff[ 731: 728] = ({4{loc_sram_buff_w0[73][4]}} & loc_sram_buff_w0[73][3:0]) | ({4{loc_sram_buff_w1[73][4]}} & loc_sram_buff_w1[73][3:0]) | ({4{loc_sram_buff_w2[73][4]}} & loc_sram_buff_w2[73][3:0]) | ({4{loc_sram_buff_w3[73][4]}} & loc_sram_buff_w3[73][3:0]) | ({4{loc_sram_buff_w4[73][4]}} & loc_sram_buff_w4[73][3:0]) | ({4{loc_sram_buff_w5[73][4]}} & loc_sram_buff_w5[73][3:0]) | ({4{loc_sram_buff_w6[73][4]}} & loc_sram_buff_w6[73][3:0]) | ({4{loc_sram_buff_w7[73][4]}} & loc_sram_buff_w7[73][3:0]) | ({4{loc_sram_buff_w8[73][4]}} & loc_sram_buff_w8[73][3:0]) | ({4{loc_sram_buff_w9[73][4]}} & loc_sram_buff_w9[73][3:0]) | ({4{loc_sram_buff_w10[73][4]}} & loc_sram_buff_w10[73][3:0]) | ({4{loc_sram_buff_w11[73][4]}} & loc_sram_buff_w11[73][3:0]) | ({4{loc_sram_buff_w12[73][4]}} & loc_sram_buff_w12[73][3:0]) | ({4{loc_sram_buff_w13[73][4]}} & loc_sram_buff_w13[73][3:0]) | ({4{loc_sram_buff_w14[73][4]}} & loc_sram_buff_w14[73][3:0]) | ({4{loc_sram_buff_w15[73][4]}} & loc_sram_buff_w15[73][3:0]);
	loc_rdata_buff[ 727: 724] = ({4{loc_sram_buff_w0[74][4]}} & loc_sram_buff_w0[74][3:0]) | ({4{loc_sram_buff_w1[74][4]}} & loc_sram_buff_w1[74][3:0]) | ({4{loc_sram_buff_w2[74][4]}} & loc_sram_buff_w2[74][3:0]) | ({4{loc_sram_buff_w3[74][4]}} & loc_sram_buff_w3[74][3:0]) | ({4{loc_sram_buff_w4[74][4]}} & loc_sram_buff_w4[74][3:0]) | ({4{loc_sram_buff_w5[74][4]}} & loc_sram_buff_w5[74][3:0]) | ({4{loc_sram_buff_w6[74][4]}} & loc_sram_buff_w6[74][3:0]) | ({4{loc_sram_buff_w7[74][4]}} & loc_sram_buff_w7[74][3:0]) | ({4{loc_sram_buff_w8[74][4]}} & loc_sram_buff_w8[74][3:0]) | ({4{loc_sram_buff_w9[74][4]}} & loc_sram_buff_w9[74][3:0]) | ({4{loc_sram_buff_w10[74][4]}} & loc_sram_buff_w10[74][3:0]) | ({4{loc_sram_buff_w11[74][4]}} & loc_sram_buff_w11[74][3:0]) | ({4{loc_sram_buff_w12[74][4]}} & loc_sram_buff_w12[74][3:0]) | ({4{loc_sram_buff_w13[74][4]}} & loc_sram_buff_w13[74][3:0]) | ({4{loc_sram_buff_w14[74][4]}} & loc_sram_buff_w14[74][3:0]) | ({4{loc_sram_buff_w15[74][4]}} & loc_sram_buff_w15[74][3:0]);
	loc_rdata_buff[ 723: 720] = ({4{loc_sram_buff_w0[75][4]}} & loc_sram_buff_w0[75][3:0]) | ({4{loc_sram_buff_w1[75][4]}} & loc_sram_buff_w1[75][3:0]) | ({4{loc_sram_buff_w2[75][4]}} & loc_sram_buff_w2[75][3:0]) | ({4{loc_sram_buff_w3[75][4]}} & loc_sram_buff_w3[75][3:0]) | ({4{loc_sram_buff_w4[75][4]}} & loc_sram_buff_w4[75][3:0]) | ({4{loc_sram_buff_w5[75][4]}} & loc_sram_buff_w5[75][3:0]) | ({4{loc_sram_buff_w6[75][4]}} & loc_sram_buff_w6[75][3:0]) | ({4{loc_sram_buff_w7[75][4]}} & loc_sram_buff_w7[75][3:0]) | ({4{loc_sram_buff_w8[75][4]}} & loc_sram_buff_w8[75][3:0]) | ({4{loc_sram_buff_w9[75][4]}} & loc_sram_buff_w9[75][3:0]) | ({4{loc_sram_buff_w10[75][4]}} & loc_sram_buff_w10[75][3:0]) | ({4{loc_sram_buff_w11[75][4]}} & loc_sram_buff_w11[75][3:0]) | ({4{loc_sram_buff_w12[75][4]}} & loc_sram_buff_w12[75][3:0]) | ({4{loc_sram_buff_w13[75][4]}} & loc_sram_buff_w13[75][3:0]) | ({4{loc_sram_buff_w14[75][4]}} & loc_sram_buff_w14[75][3:0]) | ({4{loc_sram_buff_w15[75][4]}} & loc_sram_buff_w15[75][3:0]);
	loc_rdata_buff[ 719: 716] = ({4{loc_sram_buff_w0[76][4]}} & loc_sram_buff_w0[76][3:0]) | ({4{loc_sram_buff_w1[76][4]}} & loc_sram_buff_w1[76][3:0]) | ({4{loc_sram_buff_w2[76][4]}} & loc_sram_buff_w2[76][3:0]) | ({4{loc_sram_buff_w3[76][4]}} & loc_sram_buff_w3[76][3:0]) | ({4{loc_sram_buff_w4[76][4]}} & loc_sram_buff_w4[76][3:0]) | ({4{loc_sram_buff_w5[76][4]}} & loc_sram_buff_w5[76][3:0]) | ({4{loc_sram_buff_w6[76][4]}} & loc_sram_buff_w6[76][3:0]) | ({4{loc_sram_buff_w7[76][4]}} & loc_sram_buff_w7[76][3:0]) | ({4{loc_sram_buff_w8[76][4]}} & loc_sram_buff_w8[76][3:0]) | ({4{loc_sram_buff_w9[76][4]}} & loc_sram_buff_w9[76][3:0]) | ({4{loc_sram_buff_w10[76][4]}} & loc_sram_buff_w10[76][3:0]) | ({4{loc_sram_buff_w11[76][4]}} & loc_sram_buff_w11[76][3:0]) | ({4{loc_sram_buff_w12[76][4]}} & loc_sram_buff_w12[76][3:0]) | ({4{loc_sram_buff_w13[76][4]}} & loc_sram_buff_w13[76][3:0]) | ({4{loc_sram_buff_w14[76][4]}} & loc_sram_buff_w14[76][3:0]) | ({4{loc_sram_buff_w15[76][4]}} & loc_sram_buff_w15[76][3:0]);
	loc_rdata_buff[ 715: 712] = ({4{loc_sram_buff_w0[77][4]}} & loc_sram_buff_w0[77][3:0]) | ({4{loc_sram_buff_w1[77][4]}} & loc_sram_buff_w1[77][3:0]) | ({4{loc_sram_buff_w2[77][4]}} & loc_sram_buff_w2[77][3:0]) | ({4{loc_sram_buff_w3[77][4]}} & loc_sram_buff_w3[77][3:0]) | ({4{loc_sram_buff_w4[77][4]}} & loc_sram_buff_w4[77][3:0]) | ({4{loc_sram_buff_w5[77][4]}} & loc_sram_buff_w5[77][3:0]) | ({4{loc_sram_buff_w6[77][4]}} & loc_sram_buff_w6[77][3:0]) | ({4{loc_sram_buff_w7[77][4]}} & loc_sram_buff_w7[77][3:0]) | ({4{loc_sram_buff_w8[77][4]}} & loc_sram_buff_w8[77][3:0]) | ({4{loc_sram_buff_w9[77][4]}} & loc_sram_buff_w9[77][3:0]) | ({4{loc_sram_buff_w10[77][4]}} & loc_sram_buff_w10[77][3:0]) | ({4{loc_sram_buff_w11[77][4]}} & loc_sram_buff_w11[77][3:0]) | ({4{loc_sram_buff_w12[77][4]}} & loc_sram_buff_w12[77][3:0]) | ({4{loc_sram_buff_w13[77][4]}} & loc_sram_buff_w13[77][3:0]) | ({4{loc_sram_buff_w14[77][4]}} & loc_sram_buff_w14[77][3:0]) | ({4{loc_sram_buff_w15[77][4]}} & loc_sram_buff_w15[77][3:0]);
	loc_rdata_buff[ 711: 708] = ({4{loc_sram_buff_w0[78][4]}} & loc_sram_buff_w0[78][3:0]) | ({4{loc_sram_buff_w1[78][4]}} & loc_sram_buff_w1[78][3:0]) | ({4{loc_sram_buff_w2[78][4]}} & loc_sram_buff_w2[78][3:0]) | ({4{loc_sram_buff_w3[78][4]}} & loc_sram_buff_w3[78][3:0]) | ({4{loc_sram_buff_w4[78][4]}} & loc_sram_buff_w4[78][3:0]) | ({4{loc_sram_buff_w5[78][4]}} & loc_sram_buff_w5[78][3:0]) | ({4{loc_sram_buff_w6[78][4]}} & loc_sram_buff_w6[78][3:0]) | ({4{loc_sram_buff_w7[78][4]}} & loc_sram_buff_w7[78][3:0]) | ({4{loc_sram_buff_w8[78][4]}} & loc_sram_buff_w8[78][3:0]) | ({4{loc_sram_buff_w9[78][4]}} & loc_sram_buff_w9[78][3:0]) | ({4{loc_sram_buff_w10[78][4]}} & loc_sram_buff_w10[78][3:0]) | ({4{loc_sram_buff_w11[78][4]}} & loc_sram_buff_w11[78][3:0]) | ({4{loc_sram_buff_w12[78][4]}} & loc_sram_buff_w12[78][3:0]) | ({4{loc_sram_buff_w13[78][4]}} & loc_sram_buff_w13[78][3:0]) | ({4{loc_sram_buff_w14[78][4]}} & loc_sram_buff_w14[78][3:0]) | ({4{loc_sram_buff_w15[78][4]}} & loc_sram_buff_w15[78][3:0]);
	loc_rdata_buff[ 707: 704] = ({4{loc_sram_buff_w0[79][4]}} & loc_sram_buff_w0[79][3:0]) | ({4{loc_sram_buff_w1[79][4]}} & loc_sram_buff_w1[79][3:0]) | ({4{loc_sram_buff_w2[79][4]}} & loc_sram_buff_w2[79][3:0]) | ({4{loc_sram_buff_w3[79][4]}} & loc_sram_buff_w3[79][3:0]) | ({4{loc_sram_buff_w4[79][4]}} & loc_sram_buff_w4[79][3:0]) | ({4{loc_sram_buff_w5[79][4]}} & loc_sram_buff_w5[79][3:0]) | ({4{loc_sram_buff_w6[79][4]}} & loc_sram_buff_w6[79][3:0]) | ({4{loc_sram_buff_w7[79][4]}} & loc_sram_buff_w7[79][3:0]) | ({4{loc_sram_buff_w8[79][4]}} & loc_sram_buff_w8[79][3:0]) | ({4{loc_sram_buff_w9[79][4]}} & loc_sram_buff_w9[79][3:0]) | ({4{loc_sram_buff_w10[79][4]}} & loc_sram_buff_w10[79][3:0]) | ({4{loc_sram_buff_w11[79][4]}} & loc_sram_buff_w11[79][3:0]) | ({4{loc_sram_buff_w12[79][4]}} & loc_sram_buff_w12[79][3:0]) | ({4{loc_sram_buff_w13[79][4]}} & loc_sram_buff_w13[79][3:0]) | ({4{loc_sram_buff_w14[79][4]}} & loc_sram_buff_w14[79][3:0]) | ({4{loc_sram_buff_w15[79][4]}} & loc_sram_buff_w15[79][3:0]);
	loc_rdata_buff[ 703: 700] = ({4{loc_sram_buff_w0[80][4]}} & loc_sram_buff_w0[80][3:0]) | ({4{loc_sram_buff_w1[80][4]}} & loc_sram_buff_w1[80][3:0]) | ({4{loc_sram_buff_w2[80][4]}} & loc_sram_buff_w2[80][3:0]) | ({4{loc_sram_buff_w3[80][4]}} & loc_sram_buff_w3[80][3:0]) | ({4{loc_sram_buff_w4[80][4]}} & loc_sram_buff_w4[80][3:0]) | ({4{loc_sram_buff_w5[80][4]}} & loc_sram_buff_w5[80][3:0]) | ({4{loc_sram_buff_w6[80][4]}} & loc_sram_buff_w6[80][3:0]) | ({4{loc_sram_buff_w7[80][4]}} & loc_sram_buff_w7[80][3:0]) | ({4{loc_sram_buff_w8[80][4]}} & loc_sram_buff_w8[80][3:0]) | ({4{loc_sram_buff_w9[80][4]}} & loc_sram_buff_w9[80][3:0]) | ({4{loc_sram_buff_w10[80][4]}} & loc_sram_buff_w10[80][3:0]) | ({4{loc_sram_buff_w11[80][4]}} & loc_sram_buff_w11[80][3:0]) | ({4{loc_sram_buff_w12[80][4]}} & loc_sram_buff_w12[80][3:0]) | ({4{loc_sram_buff_w13[80][4]}} & loc_sram_buff_w13[80][3:0]) | ({4{loc_sram_buff_w14[80][4]}} & loc_sram_buff_w14[80][3:0]) | ({4{loc_sram_buff_w15[80][4]}} & loc_sram_buff_w15[80][3:0]);
	loc_rdata_buff[ 699: 696] = ({4{loc_sram_buff_w0[81][4]}} & loc_sram_buff_w0[81][3:0]) | ({4{loc_sram_buff_w1[81][4]}} & loc_sram_buff_w1[81][3:0]) | ({4{loc_sram_buff_w2[81][4]}} & loc_sram_buff_w2[81][3:0]) | ({4{loc_sram_buff_w3[81][4]}} & loc_sram_buff_w3[81][3:0]) | ({4{loc_sram_buff_w4[81][4]}} & loc_sram_buff_w4[81][3:0]) | ({4{loc_sram_buff_w5[81][4]}} & loc_sram_buff_w5[81][3:0]) | ({4{loc_sram_buff_w6[81][4]}} & loc_sram_buff_w6[81][3:0]) | ({4{loc_sram_buff_w7[81][4]}} & loc_sram_buff_w7[81][3:0]) | ({4{loc_sram_buff_w8[81][4]}} & loc_sram_buff_w8[81][3:0]) | ({4{loc_sram_buff_w9[81][4]}} & loc_sram_buff_w9[81][3:0]) | ({4{loc_sram_buff_w10[81][4]}} & loc_sram_buff_w10[81][3:0]) | ({4{loc_sram_buff_w11[81][4]}} & loc_sram_buff_w11[81][3:0]) | ({4{loc_sram_buff_w12[81][4]}} & loc_sram_buff_w12[81][3:0]) | ({4{loc_sram_buff_w13[81][4]}} & loc_sram_buff_w13[81][3:0]) | ({4{loc_sram_buff_w14[81][4]}} & loc_sram_buff_w14[81][3:0]) | ({4{loc_sram_buff_w15[81][4]}} & loc_sram_buff_w15[81][3:0]);
	loc_rdata_buff[ 695: 692] = ({4{loc_sram_buff_w0[82][4]}} & loc_sram_buff_w0[82][3:0]) | ({4{loc_sram_buff_w1[82][4]}} & loc_sram_buff_w1[82][3:0]) | ({4{loc_sram_buff_w2[82][4]}} & loc_sram_buff_w2[82][3:0]) | ({4{loc_sram_buff_w3[82][4]}} & loc_sram_buff_w3[82][3:0]) | ({4{loc_sram_buff_w4[82][4]}} & loc_sram_buff_w4[82][3:0]) | ({4{loc_sram_buff_w5[82][4]}} & loc_sram_buff_w5[82][3:0]) | ({4{loc_sram_buff_w6[82][4]}} & loc_sram_buff_w6[82][3:0]) | ({4{loc_sram_buff_w7[82][4]}} & loc_sram_buff_w7[82][3:0]) | ({4{loc_sram_buff_w8[82][4]}} & loc_sram_buff_w8[82][3:0]) | ({4{loc_sram_buff_w9[82][4]}} & loc_sram_buff_w9[82][3:0]) | ({4{loc_sram_buff_w10[82][4]}} & loc_sram_buff_w10[82][3:0]) | ({4{loc_sram_buff_w11[82][4]}} & loc_sram_buff_w11[82][3:0]) | ({4{loc_sram_buff_w12[82][4]}} & loc_sram_buff_w12[82][3:0]) | ({4{loc_sram_buff_w13[82][4]}} & loc_sram_buff_w13[82][3:0]) | ({4{loc_sram_buff_w14[82][4]}} & loc_sram_buff_w14[82][3:0]) | ({4{loc_sram_buff_w15[82][4]}} & loc_sram_buff_w15[82][3:0]);
	loc_rdata_buff[ 691: 688] = ({4{loc_sram_buff_w0[83][4]}} & loc_sram_buff_w0[83][3:0]) | ({4{loc_sram_buff_w1[83][4]}} & loc_sram_buff_w1[83][3:0]) | ({4{loc_sram_buff_w2[83][4]}} & loc_sram_buff_w2[83][3:0]) | ({4{loc_sram_buff_w3[83][4]}} & loc_sram_buff_w3[83][3:0]) | ({4{loc_sram_buff_w4[83][4]}} & loc_sram_buff_w4[83][3:0]) | ({4{loc_sram_buff_w5[83][4]}} & loc_sram_buff_w5[83][3:0]) | ({4{loc_sram_buff_w6[83][4]}} & loc_sram_buff_w6[83][3:0]) | ({4{loc_sram_buff_w7[83][4]}} & loc_sram_buff_w7[83][3:0]) | ({4{loc_sram_buff_w8[83][4]}} & loc_sram_buff_w8[83][3:0]) | ({4{loc_sram_buff_w9[83][4]}} & loc_sram_buff_w9[83][3:0]) | ({4{loc_sram_buff_w10[83][4]}} & loc_sram_buff_w10[83][3:0]) | ({4{loc_sram_buff_w11[83][4]}} & loc_sram_buff_w11[83][3:0]) | ({4{loc_sram_buff_w12[83][4]}} & loc_sram_buff_w12[83][3:0]) | ({4{loc_sram_buff_w13[83][4]}} & loc_sram_buff_w13[83][3:0]) | ({4{loc_sram_buff_w14[83][4]}} & loc_sram_buff_w14[83][3:0]) | ({4{loc_sram_buff_w15[83][4]}} & loc_sram_buff_w15[83][3:0]);
	loc_rdata_buff[ 687: 684] = ({4{loc_sram_buff_w0[84][4]}} & loc_sram_buff_w0[84][3:0]) | ({4{loc_sram_buff_w1[84][4]}} & loc_sram_buff_w1[84][3:0]) | ({4{loc_sram_buff_w2[84][4]}} & loc_sram_buff_w2[84][3:0]) | ({4{loc_sram_buff_w3[84][4]}} & loc_sram_buff_w3[84][3:0]) | ({4{loc_sram_buff_w4[84][4]}} & loc_sram_buff_w4[84][3:0]) | ({4{loc_sram_buff_w5[84][4]}} & loc_sram_buff_w5[84][3:0]) | ({4{loc_sram_buff_w6[84][4]}} & loc_sram_buff_w6[84][3:0]) | ({4{loc_sram_buff_w7[84][4]}} & loc_sram_buff_w7[84][3:0]) | ({4{loc_sram_buff_w8[84][4]}} & loc_sram_buff_w8[84][3:0]) | ({4{loc_sram_buff_w9[84][4]}} & loc_sram_buff_w9[84][3:0]) | ({4{loc_sram_buff_w10[84][4]}} & loc_sram_buff_w10[84][3:0]) | ({4{loc_sram_buff_w11[84][4]}} & loc_sram_buff_w11[84][3:0]) | ({4{loc_sram_buff_w12[84][4]}} & loc_sram_buff_w12[84][3:0]) | ({4{loc_sram_buff_w13[84][4]}} & loc_sram_buff_w13[84][3:0]) | ({4{loc_sram_buff_w14[84][4]}} & loc_sram_buff_w14[84][3:0]) | ({4{loc_sram_buff_w15[84][4]}} & loc_sram_buff_w15[84][3:0]);
	loc_rdata_buff[ 683: 680] = ({4{loc_sram_buff_w0[85][4]}} & loc_sram_buff_w0[85][3:0]) | ({4{loc_sram_buff_w1[85][4]}} & loc_sram_buff_w1[85][3:0]) | ({4{loc_sram_buff_w2[85][4]}} & loc_sram_buff_w2[85][3:0]) | ({4{loc_sram_buff_w3[85][4]}} & loc_sram_buff_w3[85][3:0]) | ({4{loc_sram_buff_w4[85][4]}} & loc_sram_buff_w4[85][3:0]) | ({4{loc_sram_buff_w5[85][4]}} & loc_sram_buff_w5[85][3:0]) | ({4{loc_sram_buff_w6[85][4]}} & loc_sram_buff_w6[85][3:0]) | ({4{loc_sram_buff_w7[85][4]}} & loc_sram_buff_w7[85][3:0]) | ({4{loc_sram_buff_w8[85][4]}} & loc_sram_buff_w8[85][3:0]) | ({4{loc_sram_buff_w9[85][4]}} & loc_sram_buff_w9[85][3:0]) | ({4{loc_sram_buff_w10[85][4]}} & loc_sram_buff_w10[85][3:0]) | ({4{loc_sram_buff_w11[85][4]}} & loc_sram_buff_w11[85][3:0]) | ({4{loc_sram_buff_w12[85][4]}} & loc_sram_buff_w12[85][3:0]) | ({4{loc_sram_buff_w13[85][4]}} & loc_sram_buff_w13[85][3:0]) | ({4{loc_sram_buff_w14[85][4]}} & loc_sram_buff_w14[85][3:0]) | ({4{loc_sram_buff_w15[85][4]}} & loc_sram_buff_w15[85][3:0]);
	loc_rdata_buff[ 679: 676] = ({4{loc_sram_buff_w0[86][4]}} & loc_sram_buff_w0[86][3:0]) | ({4{loc_sram_buff_w1[86][4]}} & loc_sram_buff_w1[86][3:0]) | ({4{loc_sram_buff_w2[86][4]}} & loc_sram_buff_w2[86][3:0]) | ({4{loc_sram_buff_w3[86][4]}} & loc_sram_buff_w3[86][3:0]) | ({4{loc_sram_buff_w4[86][4]}} & loc_sram_buff_w4[86][3:0]) | ({4{loc_sram_buff_w5[86][4]}} & loc_sram_buff_w5[86][3:0]) | ({4{loc_sram_buff_w6[86][4]}} & loc_sram_buff_w6[86][3:0]) | ({4{loc_sram_buff_w7[86][4]}} & loc_sram_buff_w7[86][3:0]) | ({4{loc_sram_buff_w8[86][4]}} & loc_sram_buff_w8[86][3:0]) | ({4{loc_sram_buff_w9[86][4]}} & loc_sram_buff_w9[86][3:0]) | ({4{loc_sram_buff_w10[86][4]}} & loc_sram_buff_w10[86][3:0]) | ({4{loc_sram_buff_w11[86][4]}} & loc_sram_buff_w11[86][3:0]) | ({4{loc_sram_buff_w12[86][4]}} & loc_sram_buff_w12[86][3:0]) | ({4{loc_sram_buff_w13[86][4]}} & loc_sram_buff_w13[86][3:0]) | ({4{loc_sram_buff_w14[86][4]}} & loc_sram_buff_w14[86][3:0]) | ({4{loc_sram_buff_w15[86][4]}} & loc_sram_buff_w15[86][3:0]);
	loc_rdata_buff[ 675: 672] = ({4{loc_sram_buff_w0[87][4]}} & loc_sram_buff_w0[87][3:0]) | ({4{loc_sram_buff_w1[87][4]}} & loc_sram_buff_w1[87][3:0]) | ({4{loc_sram_buff_w2[87][4]}} & loc_sram_buff_w2[87][3:0]) | ({4{loc_sram_buff_w3[87][4]}} & loc_sram_buff_w3[87][3:0]) | ({4{loc_sram_buff_w4[87][4]}} & loc_sram_buff_w4[87][3:0]) | ({4{loc_sram_buff_w5[87][4]}} & loc_sram_buff_w5[87][3:0]) | ({4{loc_sram_buff_w6[87][4]}} & loc_sram_buff_w6[87][3:0]) | ({4{loc_sram_buff_w7[87][4]}} & loc_sram_buff_w7[87][3:0]) | ({4{loc_sram_buff_w8[87][4]}} & loc_sram_buff_w8[87][3:0]) | ({4{loc_sram_buff_w9[87][4]}} & loc_sram_buff_w9[87][3:0]) | ({4{loc_sram_buff_w10[87][4]}} & loc_sram_buff_w10[87][3:0]) | ({4{loc_sram_buff_w11[87][4]}} & loc_sram_buff_w11[87][3:0]) | ({4{loc_sram_buff_w12[87][4]}} & loc_sram_buff_w12[87][3:0]) | ({4{loc_sram_buff_w13[87][4]}} & loc_sram_buff_w13[87][3:0]) | ({4{loc_sram_buff_w14[87][4]}} & loc_sram_buff_w14[87][3:0]) | ({4{loc_sram_buff_w15[87][4]}} & loc_sram_buff_w15[87][3:0]);
	loc_rdata_buff[ 671: 668] = ({4{loc_sram_buff_w0[88][4]}} & loc_sram_buff_w0[88][3:0]) | ({4{loc_sram_buff_w1[88][4]}} & loc_sram_buff_w1[88][3:0]) | ({4{loc_sram_buff_w2[88][4]}} & loc_sram_buff_w2[88][3:0]) | ({4{loc_sram_buff_w3[88][4]}} & loc_sram_buff_w3[88][3:0]) | ({4{loc_sram_buff_w4[88][4]}} & loc_sram_buff_w4[88][3:0]) | ({4{loc_sram_buff_w5[88][4]}} & loc_sram_buff_w5[88][3:0]) | ({4{loc_sram_buff_w6[88][4]}} & loc_sram_buff_w6[88][3:0]) | ({4{loc_sram_buff_w7[88][4]}} & loc_sram_buff_w7[88][3:0]) | ({4{loc_sram_buff_w8[88][4]}} & loc_sram_buff_w8[88][3:0]) | ({4{loc_sram_buff_w9[88][4]}} & loc_sram_buff_w9[88][3:0]) | ({4{loc_sram_buff_w10[88][4]}} & loc_sram_buff_w10[88][3:0]) | ({4{loc_sram_buff_w11[88][4]}} & loc_sram_buff_w11[88][3:0]) | ({4{loc_sram_buff_w12[88][4]}} & loc_sram_buff_w12[88][3:0]) | ({4{loc_sram_buff_w13[88][4]}} & loc_sram_buff_w13[88][3:0]) | ({4{loc_sram_buff_w14[88][4]}} & loc_sram_buff_w14[88][3:0]) | ({4{loc_sram_buff_w15[88][4]}} & loc_sram_buff_w15[88][3:0]);
	loc_rdata_buff[ 667: 664] = ({4{loc_sram_buff_w0[89][4]}} & loc_sram_buff_w0[89][3:0]) | ({4{loc_sram_buff_w1[89][4]}} & loc_sram_buff_w1[89][3:0]) | ({4{loc_sram_buff_w2[89][4]}} & loc_sram_buff_w2[89][3:0]) | ({4{loc_sram_buff_w3[89][4]}} & loc_sram_buff_w3[89][3:0]) | ({4{loc_sram_buff_w4[89][4]}} & loc_sram_buff_w4[89][3:0]) | ({4{loc_sram_buff_w5[89][4]}} & loc_sram_buff_w5[89][3:0]) | ({4{loc_sram_buff_w6[89][4]}} & loc_sram_buff_w6[89][3:0]) | ({4{loc_sram_buff_w7[89][4]}} & loc_sram_buff_w7[89][3:0]) | ({4{loc_sram_buff_w8[89][4]}} & loc_sram_buff_w8[89][3:0]) | ({4{loc_sram_buff_w9[89][4]}} & loc_sram_buff_w9[89][3:0]) | ({4{loc_sram_buff_w10[89][4]}} & loc_sram_buff_w10[89][3:0]) | ({4{loc_sram_buff_w11[89][4]}} & loc_sram_buff_w11[89][3:0]) | ({4{loc_sram_buff_w12[89][4]}} & loc_sram_buff_w12[89][3:0]) | ({4{loc_sram_buff_w13[89][4]}} & loc_sram_buff_w13[89][3:0]) | ({4{loc_sram_buff_w14[89][4]}} & loc_sram_buff_w14[89][3:0]) | ({4{loc_sram_buff_w15[89][4]}} & loc_sram_buff_w15[89][3:0]);
	loc_rdata_buff[ 663: 660] = ({4{loc_sram_buff_w0[90][4]}} & loc_sram_buff_w0[90][3:0]) | ({4{loc_sram_buff_w1[90][4]}} & loc_sram_buff_w1[90][3:0]) | ({4{loc_sram_buff_w2[90][4]}} & loc_sram_buff_w2[90][3:0]) | ({4{loc_sram_buff_w3[90][4]}} & loc_sram_buff_w3[90][3:0]) | ({4{loc_sram_buff_w4[90][4]}} & loc_sram_buff_w4[90][3:0]) | ({4{loc_sram_buff_w5[90][4]}} & loc_sram_buff_w5[90][3:0]) | ({4{loc_sram_buff_w6[90][4]}} & loc_sram_buff_w6[90][3:0]) | ({4{loc_sram_buff_w7[90][4]}} & loc_sram_buff_w7[90][3:0]) | ({4{loc_sram_buff_w8[90][4]}} & loc_sram_buff_w8[90][3:0]) | ({4{loc_sram_buff_w9[90][4]}} & loc_sram_buff_w9[90][3:0]) | ({4{loc_sram_buff_w10[90][4]}} & loc_sram_buff_w10[90][3:0]) | ({4{loc_sram_buff_w11[90][4]}} & loc_sram_buff_w11[90][3:0]) | ({4{loc_sram_buff_w12[90][4]}} & loc_sram_buff_w12[90][3:0]) | ({4{loc_sram_buff_w13[90][4]}} & loc_sram_buff_w13[90][3:0]) | ({4{loc_sram_buff_w14[90][4]}} & loc_sram_buff_w14[90][3:0]) | ({4{loc_sram_buff_w15[90][4]}} & loc_sram_buff_w15[90][3:0]);
	loc_rdata_buff[ 659: 656] = ({4{loc_sram_buff_w0[91][4]}} & loc_sram_buff_w0[91][3:0]) | ({4{loc_sram_buff_w1[91][4]}} & loc_sram_buff_w1[91][3:0]) | ({4{loc_sram_buff_w2[91][4]}} & loc_sram_buff_w2[91][3:0]) | ({4{loc_sram_buff_w3[91][4]}} & loc_sram_buff_w3[91][3:0]) | ({4{loc_sram_buff_w4[91][4]}} & loc_sram_buff_w4[91][3:0]) | ({4{loc_sram_buff_w5[91][4]}} & loc_sram_buff_w5[91][3:0]) | ({4{loc_sram_buff_w6[91][4]}} & loc_sram_buff_w6[91][3:0]) | ({4{loc_sram_buff_w7[91][4]}} & loc_sram_buff_w7[91][3:0]) | ({4{loc_sram_buff_w8[91][4]}} & loc_sram_buff_w8[91][3:0]) | ({4{loc_sram_buff_w9[91][4]}} & loc_sram_buff_w9[91][3:0]) | ({4{loc_sram_buff_w10[91][4]}} & loc_sram_buff_w10[91][3:0]) | ({4{loc_sram_buff_w11[91][4]}} & loc_sram_buff_w11[91][3:0]) | ({4{loc_sram_buff_w12[91][4]}} & loc_sram_buff_w12[91][3:0]) | ({4{loc_sram_buff_w13[91][4]}} & loc_sram_buff_w13[91][3:0]) | ({4{loc_sram_buff_w14[91][4]}} & loc_sram_buff_w14[91][3:0]) | ({4{loc_sram_buff_w15[91][4]}} & loc_sram_buff_w15[91][3:0]);
	loc_rdata_buff[ 655: 652] = ({4{loc_sram_buff_w0[92][4]}} & loc_sram_buff_w0[92][3:0]) | ({4{loc_sram_buff_w1[92][4]}} & loc_sram_buff_w1[92][3:0]) | ({4{loc_sram_buff_w2[92][4]}} & loc_sram_buff_w2[92][3:0]) | ({4{loc_sram_buff_w3[92][4]}} & loc_sram_buff_w3[92][3:0]) | ({4{loc_sram_buff_w4[92][4]}} & loc_sram_buff_w4[92][3:0]) | ({4{loc_sram_buff_w5[92][4]}} & loc_sram_buff_w5[92][3:0]) | ({4{loc_sram_buff_w6[92][4]}} & loc_sram_buff_w6[92][3:0]) | ({4{loc_sram_buff_w7[92][4]}} & loc_sram_buff_w7[92][3:0]) | ({4{loc_sram_buff_w8[92][4]}} & loc_sram_buff_w8[92][3:0]) | ({4{loc_sram_buff_w9[92][4]}} & loc_sram_buff_w9[92][3:0]) | ({4{loc_sram_buff_w10[92][4]}} & loc_sram_buff_w10[92][3:0]) | ({4{loc_sram_buff_w11[92][4]}} & loc_sram_buff_w11[92][3:0]) | ({4{loc_sram_buff_w12[92][4]}} & loc_sram_buff_w12[92][3:0]) | ({4{loc_sram_buff_w13[92][4]}} & loc_sram_buff_w13[92][3:0]) | ({4{loc_sram_buff_w14[92][4]}} & loc_sram_buff_w14[92][3:0]) | ({4{loc_sram_buff_w15[92][4]}} & loc_sram_buff_w15[92][3:0]);
	loc_rdata_buff[ 651: 648] = ({4{loc_sram_buff_w0[93][4]}} & loc_sram_buff_w0[93][3:0]) | ({4{loc_sram_buff_w1[93][4]}} & loc_sram_buff_w1[93][3:0]) | ({4{loc_sram_buff_w2[93][4]}} & loc_sram_buff_w2[93][3:0]) | ({4{loc_sram_buff_w3[93][4]}} & loc_sram_buff_w3[93][3:0]) | ({4{loc_sram_buff_w4[93][4]}} & loc_sram_buff_w4[93][3:0]) | ({4{loc_sram_buff_w5[93][4]}} & loc_sram_buff_w5[93][3:0]) | ({4{loc_sram_buff_w6[93][4]}} & loc_sram_buff_w6[93][3:0]) | ({4{loc_sram_buff_w7[93][4]}} & loc_sram_buff_w7[93][3:0]) | ({4{loc_sram_buff_w8[93][4]}} & loc_sram_buff_w8[93][3:0]) | ({4{loc_sram_buff_w9[93][4]}} & loc_sram_buff_w9[93][3:0]) | ({4{loc_sram_buff_w10[93][4]}} & loc_sram_buff_w10[93][3:0]) | ({4{loc_sram_buff_w11[93][4]}} & loc_sram_buff_w11[93][3:0]) | ({4{loc_sram_buff_w12[93][4]}} & loc_sram_buff_w12[93][3:0]) | ({4{loc_sram_buff_w13[93][4]}} & loc_sram_buff_w13[93][3:0]) | ({4{loc_sram_buff_w14[93][4]}} & loc_sram_buff_w14[93][3:0]) | ({4{loc_sram_buff_w15[93][4]}} & loc_sram_buff_w15[93][3:0]);
	loc_rdata_buff[ 647: 644] = ({4{loc_sram_buff_w0[94][4]}} & loc_sram_buff_w0[94][3:0]) | ({4{loc_sram_buff_w1[94][4]}} & loc_sram_buff_w1[94][3:0]) | ({4{loc_sram_buff_w2[94][4]}} & loc_sram_buff_w2[94][3:0]) | ({4{loc_sram_buff_w3[94][4]}} & loc_sram_buff_w3[94][3:0]) | ({4{loc_sram_buff_w4[94][4]}} & loc_sram_buff_w4[94][3:0]) | ({4{loc_sram_buff_w5[94][4]}} & loc_sram_buff_w5[94][3:0]) | ({4{loc_sram_buff_w6[94][4]}} & loc_sram_buff_w6[94][3:0]) | ({4{loc_sram_buff_w7[94][4]}} & loc_sram_buff_w7[94][3:0]) | ({4{loc_sram_buff_w8[94][4]}} & loc_sram_buff_w8[94][3:0]) | ({4{loc_sram_buff_w9[94][4]}} & loc_sram_buff_w9[94][3:0]) | ({4{loc_sram_buff_w10[94][4]}} & loc_sram_buff_w10[94][3:0]) | ({4{loc_sram_buff_w11[94][4]}} & loc_sram_buff_w11[94][3:0]) | ({4{loc_sram_buff_w12[94][4]}} & loc_sram_buff_w12[94][3:0]) | ({4{loc_sram_buff_w13[94][4]}} & loc_sram_buff_w13[94][3:0]) | ({4{loc_sram_buff_w14[94][4]}} & loc_sram_buff_w14[94][3:0]) | ({4{loc_sram_buff_w15[94][4]}} & loc_sram_buff_w15[94][3:0]);
	loc_rdata_buff[ 643: 640] = ({4{loc_sram_buff_w0[95][4]}} & loc_sram_buff_w0[95][3:0]) | ({4{loc_sram_buff_w1[95][4]}} & loc_sram_buff_w1[95][3:0]) | ({4{loc_sram_buff_w2[95][4]}} & loc_sram_buff_w2[95][3:0]) | ({4{loc_sram_buff_w3[95][4]}} & loc_sram_buff_w3[95][3:0]) | ({4{loc_sram_buff_w4[95][4]}} & loc_sram_buff_w4[95][3:0]) | ({4{loc_sram_buff_w5[95][4]}} & loc_sram_buff_w5[95][3:0]) | ({4{loc_sram_buff_w6[95][4]}} & loc_sram_buff_w6[95][3:0]) | ({4{loc_sram_buff_w7[95][4]}} & loc_sram_buff_w7[95][3:0]) | ({4{loc_sram_buff_w8[95][4]}} & loc_sram_buff_w8[95][3:0]) | ({4{loc_sram_buff_w9[95][4]}} & loc_sram_buff_w9[95][3:0]) | ({4{loc_sram_buff_w10[95][4]}} & loc_sram_buff_w10[95][3:0]) | ({4{loc_sram_buff_w11[95][4]}} & loc_sram_buff_w11[95][3:0]) | ({4{loc_sram_buff_w12[95][4]}} & loc_sram_buff_w12[95][3:0]) | ({4{loc_sram_buff_w13[95][4]}} & loc_sram_buff_w13[95][3:0]) | ({4{loc_sram_buff_w14[95][4]}} & loc_sram_buff_w14[95][3:0]) | ({4{loc_sram_buff_w15[95][4]}} & loc_sram_buff_w15[95][3:0]);
	loc_rdata_buff[ 639: 636] = ({4{loc_sram_buff_w0[96][4]}} & loc_sram_buff_w0[96][3:0]) | ({4{loc_sram_buff_w1[96][4]}} & loc_sram_buff_w1[96][3:0]) | ({4{loc_sram_buff_w2[96][4]}} & loc_sram_buff_w2[96][3:0]) | ({4{loc_sram_buff_w3[96][4]}} & loc_sram_buff_w3[96][3:0]) | ({4{loc_sram_buff_w4[96][4]}} & loc_sram_buff_w4[96][3:0]) | ({4{loc_sram_buff_w5[96][4]}} & loc_sram_buff_w5[96][3:0]) | ({4{loc_sram_buff_w6[96][4]}} & loc_sram_buff_w6[96][3:0]) | ({4{loc_sram_buff_w7[96][4]}} & loc_sram_buff_w7[96][3:0]) | ({4{loc_sram_buff_w8[96][4]}} & loc_sram_buff_w8[96][3:0]) | ({4{loc_sram_buff_w9[96][4]}} & loc_sram_buff_w9[96][3:0]) | ({4{loc_sram_buff_w10[96][4]}} & loc_sram_buff_w10[96][3:0]) | ({4{loc_sram_buff_w11[96][4]}} & loc_sram_buff_w11[96][3:0]) | ({4{loc_sram_buff_w12[96][4]}} & loc_sram_buff_w12[96][3:0]) | ({4{loc_sram_buff_w13[96][4]}} & loc_sram_buff_w13[96][3:0]) | ({4{loc_sram_buff_w14[96][4]}} & loc_sram_buff_w14[96][3:0]) | ({4{loc_sram_buff_w15[96][4]}} & loc_sram_buff_w15[96][3:0]);
	loc_rdata_buff[ 635: 632] = ({4{loc_sram_buff_w0[97][4]}} & loc_sram_buff_w0[97][3:0]) | ({4{loc_sram_buff_w1[97][4]}} & loc_sram_buff_w1[97][3:0]) | ({4{loc_sram_buff_w2[97][4]}} & loc_sram_buff_w2[97][3:0]) | ({4{loc_sram_buff_w3[97][4]}} & loc_sram_buff_w3[97][3:0]) | ({4{loc_sram_buff_w4[97][4]}} & loc_sram_buff_w4[97][3:0]) | ({4{loc_sram_buff_w5[97][4]}} & loc_sram_buff_w5[97][3:0]) | ({4{loc_sram_buff_w6[97][4]}} & loc_sram_buff_w6[97][3:0]) | ({4{loc_sram_buff_w7[97][4]}} & loc_sram_buff_w7[97][3:0]) | ({4{loc_sram_buff_w8[97][4]}} & loc_sram_buff_w8[97][3:0]) | ({4{loc_sram_buff_w9[97][4]}} & loc_sram_buff_w9[97][3:0]) | ({4{loc_sram_buff_w10[97][4]}} & loc_sram_buff_w10[97][3:0]) | ({4{loc_sram_buff_w11[97][4]}} & loc_sram_buff_w11[97][3:0]) | ({4{loc_sram_buff_w12[97][4]}} & loc_sram_buff_w12[97][3:0]) | ({4{loc_sram_buff_w13[97][4]}} & loc_sram_buff_w13[97][3:0]) | ({4{loc_sram_buff_w14[97][4]}} & loc_sram_buff_w14[97][3:0]) | ({4{loc_sram_buff_w15[97][4]}} & loc_sram_buff_w15[97][3:0]);
	loc_rdata_buff[ 631: 628] = ({4{loc_sram_buff_w0[98][4]}} & loc_sram_buff_w0[98][3:0]) | ({4{loc_sram_buff_w1[98][4]}} & loc_sram_buff_w1[98][3:0]) | ({4{loc_sram_buff_w2[98][4]}} & loc_sram_buff_w2[98][3:0]) | ({4{loc_sram_buff_w3[98][4]}} & loc_sram_buff_w3[98][3:0]) | ({4{loc_sram_buff_w4[98][4]}} & loc_sram_buff_w4[98][3:0]) | ({4{loc_sram_buff_w5[98][4]}} & loc_sram_buff_w5[98][3:0]) | ({4{loc_sram_buff_w6[98][4]}} & loc_sram_buff_w6[98][3:0]) | ({4{loc_sram_buff_w7[98][4]}} & loc_sram_buff_w7[98][3:0]) | ({4{loc_sram_buff_w8[98][4]}} & loc_sram_buff_w8[98][3:0]) | ({4{loc_sram_buff_w9[98][4]}} & loc_sram_buff_w9[98][3:0]) | ({4{loc_sram_buff_w10[98][4]}} & loc_sram_buff_w10[98][3:0]) | ({4{loc_sram_buff_w11[98][4]}} & loc_sram_buff_w11[98][3:0]) | ({4{loc_sram_buff_w12[98][4]}} & loc_sram_buff_w12[98][3:0]) | ({4{loc_sram_buff_w13[98][4]}} & loc_sram_buff_w13[98][3:0]) | ({4{loc_sram_buff_w14[98][4]}} & loc_sram_buff_w14[98][3:0]) | ({4{loc_sram_buff_w15[98][4]}} & loc_sram_buff_w15[98][3:0]);
	loc_rdata_buff[ 627: 624] = ({4{loc_sram_buff_w0[99][4]}} & loc_sram_buff_w0[99][3:0]) | ({4{loc_sram_buff_w1[99][4]}} & loc_sram_buff_w1[99][3:0]) | ({4{loc_sram_buff_w2[99][4]}} & loc_sram_buff_w2[99][3:0]) | ({4{loc_sram_buff_w3[99][4]}} & loc_sram_buff_w3[99][3:0]) | ({4{loc_sram_buff_w4[99][4]}} & loc_sram_buff_w4[99][3:0]) | ({4{loc_sram_buff_w5[99][4]}} & loc_sram_buff_w5[99][3:0]) | ({4{loc_sram_buff_w6[99][4]}} & loc_sram_buff_w6[99][3:0]) | ({4{loc_sram_buff_w7[99][4]}} & loc_sram_buff_w7[99][3:0]) | ({4{loc_sram_buff_w8[99][4]}} & loc_sram_buff_w8[99][3:0]) | ({4{loc_sram_buff_w9[99][4]}} & loc_sram_buff_w9[99][3:0]) | ({4{loc_sram_buff_w10[99][4]}} & loc_sram_buff_w10[99][3:0]) | ({4{loc_sram_buff_w11[99][4]}} & loc_sram_buff_w11[99][3:0]) | ({4{loc_sram_buff_w12[99][4]}} & loc_sram_buff_w12[99][3:0]) | ({4{loc_sram_buff_w13[99][4]}} & loc_sram_buff_w13[99][3:0]) | ({4{loc_sram_buff_w14[99][4]}} & loc_sram_buff_w14[99][3:0]) | ({4{loc_sram_buff_w15[99][4]}} & loc_sram_buff_w15[99][3:0]);
	loc_rdata_buff[ 623: 620] = ({4{loc_sram_buff_w0[100][4]}} & loc_sram_buff_w0[100][3:0]) | ({4{loc_sram_buff_w1[100][4]}} & loc_sram_buff_w1[100][3:0]) | ({4{loc_sram_buff_w2[100][4]}} & loc_sram_buff_w2[100][3:0]) | ({4{loc_sram_buff_w3[100][4]}} & loc_sram_buff_w3[100][3:0]) | ({4{loc_sram_buff_w4[100][4]}} & loc_sram_buff_w4[100][3:0]) | ({4{loc_sram_buff_w5[100][4]}} & loc_sram_buff_w5[100][3:0]) | ({4{loc_sram_buff_w6[100][4]}} & loc_sram_buff_w6[100][3:0]) | ({4{loc_sram_buff_w7[100][4]}} & loc_sram_buff_w7[100][3:0]) | ({4{loc_sram_buff_w8[100][4]}} & loc_sram_buff_w8[100][3:0]) | ({4{loc_sram_buff_w9[100][4]}} & loc_sram_buff_w9[100][3:0]) | ({4{loc_sram_buff_w10[100][4]}} & loc_sram_buff_w10[100][3:0]) | ({4{loc_sram_buff_w11[100][4]}} & loc_sram_buff_w11[100][3:0]) | ({4{loc_sram_buff_w12[100][4]}} & loc_sram_buff_w12[100][3:0]) | ({4{loc_sram_buff_w13[100][4]}} & loc_sram_buff_w13[100][3:0]) | ({4{loc_sram_buff_w14[100][4]}} & loc_sram_buff_w14[100][3:0]) | ({4{loc_sram_buff_w15[100][4]}} & loc_sram_buff_w15[100][3:0]);
	loc_rdata_buff[ 619: 616] = ({4{loc_sram_buff_w0[101][4]}} & loc_sram_buff_w0[101][3:0]) | ({4{loc_sram_buff_w1[101][4]}} & loc_sram_buff_w1[101][3:0]) | ({4{loc_sram_buff_w2[101][4]}} & loc_sram_buff_w2[101][3:0]) | ({4{loc_sram_buff_w3[101][4]}} & loc_sram_buff_w3[101][3:0]) | ({4{loc_sram_buff_w4[101][4]}} & loc_sram_buff_w4[101][3:0]) | ({4{loc_sram_buff_w5[101][4]}} & loc_sram_buff_w5[101][3:0]) | ({4{loc_sram_buff_w6[101][4]}} & loc_sram_buff_w6[101][3:0]) | ({4{loc_sram_buff_w7[101][4]}} & loc_sram_buff_w7[101][3:0]) | ({4{loc_sram_buff_w8[101][4]}} & loc_sram_buff_w8[101][3:0]) | ({4{loc_sram_buff_w9[101][4]}} & loc_sram_buff_w9[101][3:0]) | ({4{loc_sram_buff_w10[101][4]}} & loc_sram_buff_w10[101][3:0]) | ({4{loc_sram_buff_w11[101][4]}} & loc_sram_buff_w11[101][3:0]) | ({4{loc_sram_buff_w12[101][4]}} & loc_sram_buff_w12[101][3:0]) | ({4{loc_sram_buff_w13[101][4]}} & loc_sram_buff_w13[101][3:0]) | ({4{loc_sram_buff_w14[101][4]}} & loc_sram_buff_w14[101][3:0]) | ({4{loc_sram_buff_w15[101][4]}} & loc_sram_buff_w15[101][3:0]);
	loc_rdata_buff[ 615: 612] = ({4{loc_sram_buff_w0[102][4]}} & loc_sram_buff_w0[102][3:0]) | ({4{loc_sram_buff_w1[102][4]}} & loc_sram_buff_w1[102][3:0]) | ({4{loc_sram_buff_w2[102][4]}} & loc_sram_buff_w2[102][3:0]) | ({4{loc_sram_buff_w3[102][4]}} & loc_sram_buff_w3[102][3:0]) | ({4{loc_sram_buff_w4[102][4]}} & loc_sram_buff_w4[102][3:0]) | ({4{loc_sram_buff_w5[102][4]}} & loc_sram_buff_w5[102][3:0]) | ({4{loc_sram_buff_w6[102][4]}} & loc_sram_buff_w6[102][3:0]) | ({4{loc_sram_buff_w7[102][4]}} & loc_sram_buff_w7[102][3:0]) | ({4{loc_sram_buff_w8[102][4]}} & loc_sram_buff_w8[102][3:0]) | ({4{loc_sram_buff_w9[102][4]}} & loc_sram_buff_w9[102][3:0]) | ({4{loc_sram_buff_w10[102][4]}} & loc_sram_buff_w10[102][3:0]) | ({4{loc_sram_buff_w11[102][4]}} & loc_sram_buff_w11[102][3:0]) | ({4{loc_sram_buff_w12[102][4]}} & loc_sram_buff_w12[102][3:0]) | ({4{loc_sram_buff_w13[102][4]}} & loc_sram_buff_w13[102][3:0]) | ({4{loc_sram_buff_w14[102][4]}} & loc_sram_buff_w14[102][3:0]) | ({4{loc_sram_buff_w15[102][4]}} & loc_sram_buff_w15[102][3:0]);
	loc_rdata_buff[ 611: 608] = ({4{loc_sram_buff_w0[103][4]}} & loc_sram_buff_w0[103][3:0]) | ({4{loc_sram_buff_w1[103][4]}} & loc_sram_buff_w1[103][3:0]) | ({4{loc_sram_buff_w2[103][4]}} & loc_sram_buff_w2[103][3:0]) | ({4{loc_sram_buff_w3[103][4]}} & loc_sram_buff_w3[103][3:0]) | ({4{loc_sram_buff_w4[103][4]}} & loc_sram_buff_w4[103][3:0]) | ({4{loc_sram_buff_w5[103][4]}} & loc_sram_buff_w5[103][3:0]) | ({4{loc_sram_buff_w6[103][4]}} & loc_sram_buff_w6[103][3:0]) | ({4{loc_sram_buff_w7[103][4]}} & loc_sram_buff_w7[103][3:0]) | ({4{loc_sram_buff_w8[103][4]}} & loc_sram_buff_w8[103][3:0]) | ({4{loc_sram_buff_w9[103][4]}} & loc_sram_buff_w9[103][3:0]) | ({4{loc_sram_buff_w10[103][4]}} & loc_sram_buff_w10[103][3:0]) | ({4{loc_sram_buff_w11[103][4]}} & loc_sram_buff_w11[103][3:0]) | ({4{loc_sram_buff_w12[103][4]}} & loc_sram_buff_w12[103][3:0]) | ({4{loc_sram_buff_w13[103][4]}} & loc_sram_buff_w13[103][3:0]) | ({4{loc_sram_buff_w14[103][4]}} & loc_sram_buff_w14[103][3:0]) | ({4{loc_sram_buff_w15[103][4]}} & loc_sram_buff_w15[103][3:0]);
	loc_rdata_buff[ 607: 604] = ({4{loc_sram_buff_w0[104][4]}} & loc_sram_buff_w0[104][3:0]) | ({4{loc_sram_buff_w1[104][4]}} & loc_sram_buff_w1[104][3:0]) | ({4{loc_sram_buff_w2[104][4]}} & loc_sram_buff_w2[104][3:0]) | ({4{loc_sram_buff_w3[104][4]}} & loc_sram_buff_w3[104][3:0]) | ({4{loc_sram_buff_w4[104][4]}} & loc_sram_buff_w4[104][3:0]) | ({4{loc_sram_buff_w5[104][4]}} & loc_sram_buff_w5[104][3:0]) | ({4{loc_sram_buff_w6[104][4]}} & loc_sram_buff_w6[104][3:0]) | ({4{loc_sram_buff_w7[104][4]}} & loc_sram_buff_w7[104][3:0]) | ({4{loc_sram_buff_w8[104][4]}} & loc_sram_buff_w8[104][3:0]) | ({4{loc_sram_buff_w9[104][4]}} & loc_sram_buff_w9[104][3:0]) | ({4{loc_sram_buff_w10[104][4]}} & loc_sram_buff_w10[104][3:0]) | ({4{loc_sram_buff_w11[104][4]}} & loc_sram_buff_w11[104][3:0]) | ({4{loc_sram_buff_w12[104][4]}} & loc_sram_buff_w12[104][3:0]) | ({4{loc_sram_buff_w13[104][4]}} & loc_sram_buff_w13[104][3:0]) | ({4{loc_sram_buff_w14[104][4]}} & loc_sram_buff_w14[104][3:0]) | ({4{loc_sram_buff_w15[104][4]}} & loc_sram_buff_w15[104][3:0]);
	loc_rdata_buff[ 603: 600] = ({4{loc_sram_buff_w0[105][4]}} & loc_sram_buff_w0[105][3:0]) | ({4{loc_sram_buff_w1[105][4]}} & loc_sram_buff_w1[105][3:0]) | ({4{loc_sram_buff_w2[105][4]}} & loc_sram_buff_w2[105][3:0]) | ({4{loc_sram_buff_w3[105][4]}} & loc_sram_buff_w3[105][3:0]) | ({4{loc_sram_buff_w4[105][4]}} & loc_sram_buff_w4[105][3:0]) | ({4{loc_sram_buff_w5[105][4]}} & loc_sram_buff_w5[105][3:0]) | ({4{loc_sram_buff_w6[105][4]}} & loc_sram_buff_w6[105][3:0]) | ({4{loc_sram_buff_w7[105][4]}} & loc_sram_buff_w7[105][3:0]) | ({4{loc_sram_buff_w8[105][4]}} & loc_sram_buff_w8[105][3:0]) | ({4{loc_sram_buff_w9[105][4]}} & loc_sram_buff_w9[105][3:0]) | ({4{loc_sram_buff_w10[105][4]}} & loc_sram_buff_w10[105][3:0]) | ({4{loc_sram_buff_w11[105][4]}} & loc_sram_buff_w11[105][3:0]) | ({4{loc_sram_buff_w12[105][4]}} & loc_sram_buff_w12[105][3:0]) | ({4{loc_sram_buff_w13[105][4]}} & loc_sram_buff_w13[105][3:0]) | ({4{loc_sram_buff_w14[105][4]}} & loc_sram_buff_w14[105][3:0]) | ({4{loc_sram_buff_w15[105][4]}} & loc_sram_buff_w15[105][3:0]);
	loc_rdata_buff[ 599: 596] = ({4{loc_sram_buff_w0[106][4]}} & loc_sram_buff_w0[106][3:0]) | ({4{loc_sram_buff_w1[106][4]}} & loc_sram_buff_w1[106][3:0]) | ({4{loc_sram_buff_w2[106][4]}} & loc_sram_buff_w2[106][3:0]) | ({4{loc_sram_buff_w3[106][4]}} & loc_sram_buff_w3[106][3:0]) | ({4{loc_sram_buff_w4[106][4]}} & loc_sram_buff_w4[106][3:0]) | ({4{loc_sram_buff_w5[106][4]}} & loc_sram_buff_w5[106][3:0]) | ({4{loc_sram_buff_w6[106][4]}} & loc_sram_buff_w6[106][3:0]) | ({4{loc_sram_buff_w7[106][4]}} & loc_sram_buff_w7[106][3:0]) | ({4{loc_sram_buff_w8[106][4]}} & loc_sram_buff_w8[106][3:0]) | ({4{loc_sram_buff_w9[106][4]}} & loc_sram_buff_w9[106][3:0]) | ({4{loc_sram_buff_w10[106][4]}} & loc_sram_buff_w10[106][3:0]) | ({4{loc_sram_buff_w11[106][4]}} & loc_sram_buff_w11[106][3:0]) | ({4{loc_sram_buff_w12[106][4]}} & loc_sram_buff_w12[106][3:0]) | ({4{loc_sram_buff_w13[106][4]}} & loc_sram_buff_w13[106][3:0]) | ({4{loc_sram_buff_w14[106][4]}} & loc_sram_buff_w14[106][3:0]) | ({4{loc_sram_buff_w15[106][4]}} & loc_sram_buff_w15[106][3:0]);
	loc_rdata_buff[ 595: 592] = ({4{loc_sram_buff_w0[107][4]}} & loc_sram_buff_w0[107][3:0]) | ({4{loc_sram_buff_w1[107][4]}} & loc_sram_buff_w1[107][3:0]) | ({4{loc_sram_buff_w2[107][4]}} & loc_sram_buff_w2[107][3:0]) | ({4{loc_sram_buff_w3[107][4]}} & loc_sram_buff_w3[107][3:0]) | ({4{loc_sram_buff_w4[107][4]}} & loc_sram_buff_w4[107][3:0]) | ({4{loc_sram_buff_w5[107][4]}} & loc_sram_buff_w5[107][3:0]) | ({4{loc_sram_buff_w6[107][4]}} & loc_sram_buff_w6[107][3:0]) | ({4{loc_sram_buff_w7[107][4]}} & loc_sram_buff_w7[107][3:0]) | ({4{loc_sram_buff_w8[107][4]}} & loc_sram_buff_w8[107][3:0]) | ({4{loc_sram_buff_w9[107][4]}} & loc_sram_buff_w9[107][3:0]) | ({4{loc_sram_buff_w10[107][4]}} & loc_sram_buff_w10[107][3:0]) | ({4{loc_sram_buff_w11[107][4]}} & loc_sram_buff_w11[107][3:0]) | ({4{loc_sram_buff_w12[107][4]}} & loc_sram_buff_w12[107][3:0]) | ({4{loc_sram_buff_w13[107][4]}} & loc_sram_buff_w13[107][3:0]) | ({4{loc_sram_buff_w14[107][4]}} & loc_sram_buff_w14[107][3:0]) | ({4{loc_sram_buff_w15[107][4]}} & loc_sram_buff_w15[107][3:0]);
	loc_rdata_buff[ 591: 588] = ({4{loc_sram_buff_w0[108][4]}} & loc_sram_buff_w0[108][3:0]) | ({4{loc_sram_buff_w1[108][4]}} & loc_sram_buff_w1[108][3:0]) | ({4{loc_sram_buff_w2[108][4]}} & loc_sram_buff_w2[108][3:0]) | ({4{loc_sram_buff_w3[108][4]}} & loc_sram_buff_w3[108][3:0]) | ({4{loc_sram_buff_w4[108][4]}} & loc_sram_buff_w4[108][3:0]) | ({4{loc_sram_buff_w5[108][4]}} & loc_sram_buff_w5[108][3:0]) | ({4{loc_sram_buff_w6[108][4]}} & loc_sram_buff_w6[108][3:0]) | ({4{loc_sram_buff_w7[108][4]}} & loc_sram_buff_w7[108][3:0]) | ({4{loc_sram_buff_w8[108][4]}} & loc_sram_buff_w8[108][3:0]) | ({4{loc_sram_buff_w9[108][4]}} & loc_sram_buff_w9[108][3:0]) | ({4{loc_sram_buff_w10[108][4]}} & loc_sram_buff_w10[108][3:0]) | ({4{loc_sram_buff_w11[108][4]}} & loc_sram_buff_w11[108][3:0]) | ({4{loc_sram_buff_w12[108][4]}} & loc_sram_buff_w12[108][3:0]) | ({4{loc_sram_buff_w13[108][4]}} & loc_sram_buff_w13[108][3:0]) | ({4{loc_sram_buff_w14[108][4]}} & loc_sram_buff_w14[108][3:0]) | ({4{loc_sram_buff_w15[108][4]}} & loc_sram_buff_w15[108][3:0]);
	loc_rdata_buff[ 587: 584] = ({4{loc_sram_buff_w0[109][4]}} & loc_sram_buff_w0[109][3:0]) | ({4{loc_sram_buff_w1[109][4]}} & loc_sram_buff_w1[109][3:0]) | ({4{loc_sram_buff_w2[109][4]}} & loc_sram_buff_w2[109][3:0]) | ({4{loc_sram_buff_w3[109][4]}} & loc_sram_buff_w3[109][3:0]) | ({4{loc_sram_buff_w4[109][4]}} & loc_sram_buff_w4[109][3:0]) | ({4{loc_sram_buff_w5[109][4]}} & loc_sram_buff_w5[109][3:0]) | ({4{loc_sram_buff_w6[109][4]}} & loc_sram_buff_w6[109][3:0]) | ({4{loc_sram_buff_w7[109][4]}} & loc_sram_buff_w7[109][3:0]) | ({4{loc_sram_buff_w8[109][4]}} & loc_sram_buff_w8[109][3:0]) | ({4{loc_sram_buff_w9[109][4]}} & loc_sram_buff_w9[109][3:0]) | ({4{loc_sram_buff_w10[109][4]}} & loc_sram_buff_w10[109][3:0]) | ({4{loc_sram_buff_w11[109][4]}} & loc_sram_buff_w11[109][3:0]) | ({4{loc_sram_buff_w12[109][4]}} & loc_sram_buff_w12[109][3:0]) | ({4{loc_sram_buff_w13[109][4]}} & loc_sram_buff_w13[109][3:0]) | ({4{loc_sram_buff_w14[109][4]}} & loc_sram_buff_w14[109][3:0]) | ({4{loc_sram_buff_w15[109][4]}} & loc_sram_buff_w15[109][3:0]);
	loc_rdata_buff[ 583: 580] = ({4{loc_sram_buff_w0[110][4]}} & loc_sram_buff_w0[110][3:0]) | ({4{loc_sram_buff_w1[110][4]}} & loc_sram_buff_w1[110][3:0]) | ({4{loc_sram_buff_w2[110][4]}} & loc_sram_buff_w2[110][3:0]) | ({4{loc_sram_buff_w3[110][4]}} & loc_sram_buff_w3[110][3:0]) | ({4{loc_sram_buff_w4[110][4]}} & loc_sram_buff_w4[110][3:0]) | ({4{loc_sram_buff_w5[110][4]}} & loc_sram_buff_w5[110][3:0]) | ({4{loc_sram_buff_w6[110][4]}} & loc_sram_buff_w6[110][3:0]) | ({4{loc_sram_buff_w7[110][4]}} & loc_sram_buff_w7[110][3:0]) | ({4{loc_sram_buff_w8[110][4]}} & loc_sram_buff_w8[110][3:0]) | ({4{loc_sram_buff_w9[110][4]}} & loc_sram_buff_w9[110][3:0]) | ({4{loc_sram_buff_w10[110][4]}} & loc_sram_buff_w10[110][3:0]) | ({4{loc_sram_buff_w11[110][4]}} & loc_sram_buff_w11[110][3:0]) | ({4{loc_sram_buff_w12[110][4]}} & loc_sram_buff_w12[110][3:0]) | ({4{loc_sram_buff_w13[110][4]}} & loc_sram_buff_w13[110][3:0]) | ({4{loc_sram_buff_w14[110][4]}} & loc_sram_buff_w14[110][3:0]) | ({4{loc_sram_buff_w15[110][4]}} & loc_sram_buff_w15[110][3:0]);
	loc_rdata_buff[ 579: 576] = ({4{loc_sram_buff_w0[111][4]}} & loc_sram_buff_w0[111][3:0]) | ({4{loc_sram_buff_w1[111][4]}} & loc_sram_buff_w1[111][3:0]) | ({4{loc_sram_buff_w2[111][4]}} & loc_sram_buff_w2[111][3:0]) | ({4{loc_sram_buff_w3[111][4]}} & loc_sram_buff_w3[111][3:0]) | ({4{loc_sram_buff_w4[111][4]}} & loc_sram_buff_w4[111][3:0]) | ({4{loc_sram_buff_w5[111][4]}} & loc_sram_buff_w5[111][3:0]) | ({4{loc_sram_buff_w6[111][4]}} & loc_sram_buff_w6[111][3:0]) | ({4{loc_sram_buff_w7[111][4]}} & loc_sram_buff_w7[111][3:0]) | ({4{loc_sram_buff_w8[111][4]}} & loc_sram_buff_w8[111][3:0]) | ({4{loc_sram_buff_w9[111][4]}} & loc_sram_buff_w9[111][3:0]) | ({4{loc_sram_buff_w10[111][4]}} & loc_sram_buff_w10[111][3:0]) | ({4{loc_sram_buff_w11[111][4]}} & loc_sram_buff_w11[111][3:0]) | ({4{loc_sram_buff_w12[111][4]}} & loc_sram_buff_w12[111][3:0]) | ({4{loc_sram_buff_w13[111][4]}} & loc_sram_buff_w13[111][3:0]) | ({4{loc_sram_buff_w14[111][4]}} & loc_sram_buff_w14[111][3:0]) | ({4{loc_sram_buff_w15[111][4]}} & loc_sram_buff_w15[111][3:0]);
	loc_rdata_buff[ 575: 572] = ({4{loc_sram_buff_w0[112][4]}} & loc_sram_buff_w0[112][3:0]) | ({4{loc_sram_buff_w1[112][4]}} & loc_sram_buff_w1[112][3:0]) | ({4{loc_sram_buff_w2[112][4]}} & loc_sram_buff_w2[112][3:0]) | ({4{loc_sram_buff_w3[112][4]}} & loc_sram_buff_w3[112][3:0]) | ({4{loc_sram_buff_w4[112][4]}} & loc_sram_buff_w4[112][3:0]) | ({4{loc_sram_buff_w5[112][4]}} & loc_sram_buff_w5[112][3:0]) | ({4{loc_sram_buff_w6[112][4]}} & loc_sram_buff_w6[112][3:0]) | ({4{loc_sram_buff_w7[112][4]}} & loc_sram_buff_w7[112][3:0]) | ({4{loc_sram_buff_w8[112][4]}} & loc_sram_buff_w8[112][3:0]) | ({4{loc_sram_buff_w9[112][4]}} & loc_sram_buff_w9[112][3:0]) | ({4{loc_sram_buff_w10[112][4]}} & loc_sram_buff_w10[112][3:0]) | ({4{loc_sram_buff_w11[112][4]}} & loc_sram_buff_w11[112][3:0]) | ({4{loc_sram_buff_w12[112][4]}} & loc_sram_buff_w12[112][3:0]) | ({4{loc_sram_buff_w13[112][4]}} & loc_sram_buff_w13[112][3:0]) | ({4{loc_sram_buff_w14[112][4]}} & loc_sram_buff_w14[112][3:0]) | ({4{loc_sram_buff_w15[112][4]}} & loc_sram_buff_w15[112][3:0]);
	loc_rdata_buff[ 571: 568] = ({4{loc_sram_buff_w0[113][4]}} & loc_sram_buff_w0[113][3:0]) | ({4{loc_sram_buff_w1[113][4]}} & loc_sram_buff_w1[113][3:0]) | ({4{loc_sram_buff_w2[113][4]}} & loc_sram_buff_w2[113][3:0]) | ({4{loc_sram_buff_w3[113][4]}} & loc_sram_buff_w3[113][3:0]) | ({4{loc_sram_buff_w4[113][4]}} & loc_sram_buff_w4[113][3:0]) | ({4{loc_sram_buff_w5[113][4]}} & loc_sram_buff_w5[113][3:0]) | ({4{loc_sram_buff_w6[113][4]}} & loc_sram_buff_w6[113][3:0]) | ({4{loc_sram_buff_w7[113][4]}} & loc_sram_buff_w7[113][3:0]) | ({4{loc_sram_buff_w8[113][4]}} & loc_sram_buff_w8[113][3:0]) | ({4{loc_sram_buff_w9[113][4]}} & loc_sram_buff_w9[113][3:0]) | ({4{loc_sram_buff_w10[113][4]}} & loc_sram_buff_w10[113][3:0]) | ({4{loc_sram_buff_w11[113][4]}} & loc_sram_buff_w11[113][3:0]) | ({4{loc_sram_buff_w12[113][4]}} & loc_sram_buff_w12[113][3:0]) | ({4{loc_sram_buff_w13[113][4]}} & loc_sram_buff_w13[113][3:0]) | ({4{loc_sram_buff_w14[113][4]}} & loc_sram_buff_w14[113][3:0]) | ({4{loc_sram_buff_w15[113][4]}} & loc_sram_buff_w15[113][3:0]);
	loc_rdata_buff[ 567: 564] = ({4{loc_sram_buff_w0[114][4]}} & loc_sram_buff_w0[114][3:0]) | ({4{loc_sram_buff_w1[114][4]}} & loc_sram_buff_w1[114][3:0]) | ({4{loc_sram_buff_w2[114][4]}} & loc_sram_buff_w2[114][3:0]) | ({4{loc_sram_buff_w3[114][4]}} & loc_sram_buff_w3[114][3:0]) | ({4{loc_sram_buff_w4[114][4]}} & loc_sram_buff_w4[114][3:0]) | ({4{loc_sram_buff_w5[114][4]}} & loc_sram_buff_w5[114][3:0]) | ({4{loc_sram_buff_w6[114][4]}} & loc_sram_buff_w6[114][3:0]) | ({4{loc_sram_buff_w7[114][4]}} & loc_sram_buff_w7[114][3:0]) | ({4{loc_sram_buff_w8[114][4]}} & loc_sram_buff_w8[114][3:0]) | ({4{loc_sram_buff_w9[114][4]}} & loc_sram_buff_w9[114][3:0]) | ({4{loc_sram_buff_w10[114][4]}} & loc_sram_buff_w10[114][3:0]) | ({4{loc_sram_buff_w11[114][4]}} & loc_sram_buff_w11[114][3:0]) | ({4{loc_sram_buff_w12[114][4]}} & loc_sram_buff_w12[114][3:0]) | ({4{loc_sram_buff_w13[114][4]}} & loc_sram_buff_w13[114][3:0]) | ({4{loc_sram_buff_w14[114][4]}} & loc_sram_buff_w14[114][3:0]) | ({4{loc_sram_buff_w15[114][4]}} & loc_sram_buff_w15[114][3:0]);
	loc_rdata_buff[ 563: 560] = ({4{loc_sram_buff_w0[115][4]}} & loc_sram_buff_w0[115][3:0]) | ({4{loc_sram_buff_w1[115][4]}} & loc_sram_buff_w1[115][3:0]) | ({4{loc_sram_buff_w2[115][4]}} & loc_sram_buff_w2[115][3:0]) | ({4{loc_sram_buff_w3[115][4]}} & loc_sram_buff_w3[115][3:0]) | ({4{loc_sram_buff_w4[115][4]}} & loc_sram_buff_w4[115][3:0]) | ({4{loc_sram_buff_w5[115][4]}} & loc_sram_buff_w5[115][3:0]) | ({4{loc_sram_buff_w6[115][4]}} & loc_sram_buff_w6[115][3:0]) | ({4{loc_sram_buff_w7[115][4]}} & loc_sram_buff_w7[115][3:0]) | ({4{loc_sram_buff_w8[115][4]}} & loc_sram_buff_w8[115][3:0]) | ({4{loc_sram_buff_w9[115][4]}} & loc_sram_buff_w9[115][3:0]) | ({4{loc_sram_buff_w10[115][4]}} & loc_sram_buff_w10[115][3:0]) | ({4{loc_sram_buff_w11[115][4]}} & loc_sram_buff_w11[115][3:0]) | ({4{loc_sram_buff_w12[115][4]}} & loc_sram_buff_w12[115][3:0]) | ({4{loc_sram_buff_w13[115][4]}} & loc_sram_buff_w13[115][3:0]) | ({4{loc_sram_buff_w14[115][4]}} & loc_sram_buff_w14[115][3:0]) | ({4{loc_sram_buff_w15[115][4]}} & loc_sram_buff_w15[115][3:0]);
	loc_rdata_buff[ 559: 556] = ({4{loc_sram_buff_w0[116][4]}} & loc_sram_buff_w0[116][3:0]) | ({4{loc_sram_buff_w1[116][4]}} & loc_sram_buff_w1[116][3:0]) | ({4{loc_sram_buff_w2[116][4]}} & loc_sram_buff_w2[116][3:0]) | ({4{loc_sram_buff_w3[116][4]}} & loc_sram_buff_w3[116][3:0]) | ({4{loc_sram_buff_w4[116][4]}} & loc_sram_buff_w4[116][3:0]) | ({4{loc_sram_buff_w5[116][4]}} & loc_sram_buff_w5[116][3:0]) | ({4{loc_sram_buff_w6[116][4]}} & loc_sram_buff_w6[116][3:0]) | ({4{loc_sram_buff_w7[116][4]}} & loc_sram_buff_w7[116][3:0]) | ({4{loc_sram_buff_w8[116][4]}} & loc_sram_buff_w8[116][3:0]) | ({4{loc_sram_buff_w9[116][4]}} & loc_sram_buff_w9[116][3:0]) | ({4{loc_sram_buff_w10[116][4]}} & loc_sram_buff_w10[116][3:0]) | ({4{loc_sram_buff_w11[116][4]}} & loc_sram_buff_w11[116][3:0]) | ({4{loc_sram_buff_w12[116][4]}} & loc_sram_buff_w12[116][3:0]) | ({4{loc_sram_buff_w13[116][4]}} & loc_sram_buff_w13[116][3:0]) | ({4{loc_sram_buff_w14[116][4]}} & loc_sram_buff_w14[116][3:0]) | ({4{loc_sram_buff_w15[116][4]}} & loc_sram_buff_w15[116][3:0]);
	loc_rdata_buff[ 555: 552] = ({4{loc_sram_buff_w0[117][4]}} & loc_sram_buff_w0[117][3:0]) | ({4{loc_sram_buff_w1[117][4]}} & loc_sram_buff_w1[117][3:0]) | ({4{loc_sram_buff_w2[117][4]}} & loc_sram_buff_w2[117][3:0]) | ({4{loc_sram_buff_w3[117][4]}} & loc_sram_buff_w3[117][3:0]) | ({4{loc_sram_buff_w4[117][4]}} & loc_sram_buff_w4[117][3:0]) | ({4{loc_sram_buff_w5[117][4]}} & loc_sram_buff_w5[117][3:0]) | ({4{loc_sram_buff_w6[117][4]}} & loc_sram_buff_w6[117][3:0]) | ({4{loc_sram_buff_w7[117][4]}} & loc_sram_buff_w7[117][3:0]) | ({4{loc_sram_buff_w8[117][4]}} & loc_sram_buff_w8[117][3:0]) | ({4{loc_sram_buff_w9[117][4]}} & loc_sram_buff_w9[117][3:0]) | ({4{loc_sram_buff_w10[117][4]}} & loc_sram_buff_w10[117][3:0]) | ({4{loc_sram_buff_w11[117][4]}} & loc_sram_buff_w11[117][3:0]) | ({4{loc_sram_buff_w12[117][4]}} & loc_sram_buff_w12[117][3:0]) | ({4{loc_sram_buff_w13[117][4]}} & loc_sram_buff_w13[117][3:0]) | ({4{loc_sram_buff_w14[117][4]}} & loc_sram_buff_w14[117][3:0]) | ({4{loc_sram_buff_w15[117][4]}} & loc_sram_buff_w15[117][3:0]);
	loc_rdata_buff[ 551: 548] = ({4{loc_sram_buff_w0[118][4]}} & loc_sram_buff_w0[118][3:0]) | ({4{loc_sram_buff_w1[118][4]}} & loc_sram_buff_w1[118][3:0]) | ({4{loc_sram_buff_w2[118][4]}} & loc_sram_buff_w2[118][3:0]) | ({4{loc_sram_buff_w3[118][4]}} & loc_sram_buff_w3[118][3:0]) | ({4{loc_sram_buff_w4[118][4]}} & loc_sram_buff_w4[118][3:0]) | ({4{loc_sram_buff_w5[118][4]}} & loc_sram_buff_w5[118][3:0]) | ({4{loc_sram_buff_w6[118][4]}} & loc_sram_buff_w6[118][3:0]) | ({4{loc_sram_buff_w7[118][4]}} & loc_sram_buff_w7[118][3:0]) | ({4{loc_sram_buff_w8[118][4]}} & loc_sram_buff_w8[118][3:0]) | ({4{loc_sram_buff_w9[118][4]}} & loc_sram_buff_w9[118][3:0]) | ({4{loc_sram_buff_w10[118][4]}} & loc_sram_buff_w10[118][3:0]) | ({4{loc_sram_buff_w11[118][4]}} & loc_sram_buff_w11[118][3:0]) | ({4{loc_sram_buff_w12[118][4]}} & loc_sram_buff_w12[118][3:0]) | ({4{loc_sram_buff_w13[118][4]}} & loc_sram_buff_w13[118][3:0]) | ({4{loc_sram_buff_w14[118][4]}} & loc_sram_buff_w14[118][3:0]) | ({4{loc_sram_buff_w15[118][4]}} & loc_sram_buff_w15[118][3:0]);
	loc_rdata_buff[ 547: 544] = ({4{loc_sram_buff_w0[119][4]}} & loc_sram_buff_w0[119][3:0]) | ({4{loc_sram_buff_w1[119][4]}} & loc_sram_buff_w1[119][3:0]) | ({4{loc_sram_buff_w2[119][4]}} & loc_sram_buff_w2[119][3:0]) | ({4{loc_sram_buff_w3[119][4]}} & loc_sram_buff_w3[119][3:0]) | ({4{loc_sram_buff_w4[119][4]}} & loc_sram_buff_w4[119][3:0]) | ({4{loc_sram_buff_w5[119][4]}} & loc_sram_buff_w5[119][3:0]) | ({4{loc_sram_buff_w6[119][4]}} & loc_sram_buff_w6[119][3:0]) | ({4{loc_sram_buff_w7[119][4]}} & loc_sram_buff_w7[119][3:0]) | ({4{loc_sram_buff_w8[119][4]}} & loc_sram_buff_w8[119][3:0]) | ({4{loc_sram_buff_w9[119][4]}} & loc_sram_buff_w9[119][3:0]) | ({4{loc_sram_buff_w10[119][4]}} & loc_sram_buff_w10[119][3:0]) | ({4{loc_sram_buff_w11[119][4]}} & loc_sram_buff_w11[119][3:0]) | ({4{loc_sram_buff_w12[119][4]}} & loc_sram_buff_w12[119][3:0]) | ({4{loc_sram_buff_w13[119][4]}} & loc_sram_buff_w13[119][3:0]) | ({4{loc_sram_buff_w14[119][4]}} & loc_sram_buff_w14[119][3:0]) | ({4{loc_sram_buff_w15[119][4]}} & loc_sram_buff_w15[119][3:0]);
	loc_rdata_buff[ 543: 540] = ({4{loc_sram_buff_w0[120][4]}} & loc_sram_buff_w0[120][3:0]) | ({4{loc_sram_buff_w1[120][4]}} & loc_sram_buff_w1[120][3:0]) | ({4{loc_sram_buff_w2[120][4]}} & loc_sram_buff_w2[120][3:0]) | ({4{loc_sram_buff_w3[120][4]}} & loc_sram_buff_w3[120][3:0]) | ({4{loc_sram_buff_w4[120][4]}} & loc_sram_buff_w4[120][3:0]) | ({4{loc_sram_buff_w5[120][4]}} & loc_sram_buff_w5[120][3:0]) | ({4{loc_sram_buff_w6[120][4]}} & loc_sram_buff_w6[120][3:0]) | ({4{loc_sram_buff_w7[120][4]}} & loc_sram_buff_w7[120][3:0]) | ({4{loc_sram_buff_w8[120][4]}} & loc_sram_buff_w8[120][3:0]) | ({4{loc_sram_buff_w9[120][4]}} & loc_sram_buff_w9[120][3:0]) | ({4{loc_sram_buff_w10[120][4]}} & loc_sram_buff_w10[120][3:0]) | ({4{loc_sram_buff_w11[120][4]}} & loc_sram_buff_w11[120][3:0]) | ({4{loc_sram_buff_w12[120][4]}} & loc_sram_buff_w12[120][3:0]) | ({4{loc_sram_buff_w13[120][4]}} & loc_sram_buff_w13[120][3:0]) | ({4{loc_sram_buff_w14[120][4]}} & loc_sram_buff_w14[120][3:0]) | ({4{loc_sram_buff_w15[120][4]}} & loc_sram_buff_w15[120][3:0]);
	loc_rdata_buff[ 539: 536] = ({4{loc_sram_buff_w0[121][4]}} & loc_sram_buff_w0[121][3:0]) | ({4{loc_sram_buff_w1[121][4]}} & loc_sram_buff_w1[121][3:0]) | ({4{loc_sram_buff_w2[121][4]}} & loc_sram_buff_w2[121][3:0]) | ({4{loc_sram_buff_w3[121][4]}} & loc_sram_buff_w3[121][3:0]) | ({4{loc_sram_buff_w4[121][4]}} & loc_sram_buff_w4[121][3:0]) | ({4{loc_sram_buff_w5[121][4]}} & loc_sram_buff_w5[121][3:0]) | ({4{loc_sram_buff_w6[121][4]}} & loc_sram_buff_w6[121][3:0]) | ({4{loc_sram_buff_w7[121][4]}} & loc_sram_buff_w7[121][3:0]) | ({4{loc_sram_buff_w8[121][4]}} & loc_sram_buff_w8[121][3:0]) | ({4{loc_sram_buff_w9[121][4]}} & loc_sram_buff_w9[121][3:0]) | ({4{loc_sram_buff_w10[121][4]}} & loc_sram_buff_w10[121][3:0]) | ({4{loc_sram_buff_w11[121][4]}} & loc_sram_buff_w11[121][3:0]) | ({4{loc_sram_buff_w12[121][4]}} & loc_sram_buff_w12[121][3:0]) | ({4{loc_sram_buff_w13[121][4]}} & loc_sram_buff_w13[121][3:0]) | ({4{loc_sram_buff_w14[121][4]}} & loc_sram_buff_w14[121][3:0]) | ({4{loc_sram_buff_w15[121][4]}} & loc_sram_buff_w15[121][3:0]);
	loc_rdata_buff[ 535: 532] = ({4{loc_sram_buff_w0[122][4]}} & loc_sram_buff_w0[122][3:0]) | ({4{loc_sram_buff_w1[122][4]}} & loc_sram_buff_w1[122][3:0]) | ({4{loc_sram_buff_w2[122][4]}} & loc_sram_buff_w2[122][3:0]) | ({4{loc_sram_buff_w3[122][4]}} & loc_sram_buff_w3[122][3:0]) | ({4{loc_sram_buff_w4[122][4]}} & loc_sram_buff_w4[122][3:0]) | ({4{loc_sram_buff_w5[122][4]}} & loc_sram_buff_w5[122][3:0]) | ({4{loc_sram_buff_w6[122][4]}} & loc_sram_buff_w6[122][3:0]) | ({4{loc_sram_buff_w7[122][4]}} & loc_sram_buff_w7[122][3:0]) | ({4{loc_sram_buff_w8[122][4]}} & loc_sram_buff_w8[122][3:0]) | ({4{loc_sram_buff_w9[122][4]}} & loc_sram_buff_w9[122][3:0]) | ({4{loc_sram_buff_w10[122][4]}} & loc_sram_buff_w10[122][3:0]) | ({4{loc_sram_buff_w11[122][4]}} & loc_sram_buff_w11[122][3:0]) | ({4{loc_sram_buff_w12[122][4]}} & loc_sram_buff_w12[122][3:0]) | ({4{loc_sram_buff_w13[122][4]}} & loc_sram_buff_w13[122][3:0]) | ({4{loc_sram_buff_w14[122][4]}} & loc_sram_buff_w14[122][3:0]) | ({4{loc_sram_buff_w15[122][4]}} & loc_sram_buff_w15[122][3:0]);
	loc_rdata_buff[ 531: 528] = ({4{loc_sram_buff_w0[123][4]}} & loc_sram_buff_w0[123][3:0]) | ({4{loc_sram_buff_w1[123][4]}} & loc_sram_buff_w1[123][3:0]) | ({4{loc_sram_buff_w2[123][4]}} & loc_sram_buff_w2[123][3:0]) | ({4{loc_sram_buff_w3[123][4]}} & loc_sram_buff_w3[123][3:0]) | ({4{loc_sram_buff_w4[123][4]}} & loc_sram_buff_w4[123][3:0]) | ({4{loc_sram_buff_w5[123][4]}} & loc_sram_buff_w5[123][3:0]) | ({4{loc_sram_buff_w6[123][4]}} & loc_sram_buff_w6[123][3:0]) | ({4{loc_sram_buff_w7[123][4]}} & loc_sram_buff_w7[123][3:0]) | ({4{loc_sram_buff_w8[123][4]}} & loc_sram_buff_w8[123][3:0]) | ({4{loc_sram_buff_w9[123][4]}} & loc_sram_buff_w9[123][3:0]) | ({4{loc_sram_buff_w10[123][4]}} & loc_sram_buff_w10[123][3:0]) | ({4{loc_sram_buff_w11[123][4]}} & loc_sram_buff_w11[123][3:0]) | ({4{loc_sram_buff_w12[123][4]}} & loc_sram_buff_w12[123][3:0]) | ({4{loc_sram_buff_w13[123][4]}} & loc_sram_buff_w13[123][3:0]) | ({4{loc_sram_buff_w14[123][4]}} & loc_sram_buff_w14[123][3:0]) | ({4{loc_sram_buff_w15[123][4]}} & loc_sram_buff_w15[123][3:0]);
	loc_rdata_buff[ 527: 524] = ({4{loc_sram_buff_w0[124][4]}} & loc_sram_buff_w0[124][3:0]) | ({4{loc_sram_buff_w1[124][4]}} & loc_sram_buff_w1[124][3:0]) | ({4{loc_sram_buff_w2[124][4]}} & loc_sram_buff_w2[124][3:0]) | ({4{loc_sram_buff_w3[124][4]}} & loc_sram_buff_w3[124][3:0]) | ({4{loc_sram_buff_w4[124][4]}} & loc_sram_buff_w4[124][3:0]) | ({4{loc_sram_buff_w5[124][4]}} & loc_sram_buff_w5[124][3:0]) | ({4{loc_sram_buff_w6[124][4]}} & loc_sram_buff_w6[124][3:0]) | ({4{loc_sram_buff_w7[124][4]}} & loc_sram_buff_w7[124][3:0]) | ({4{loc_sram_buff_w8[124][4]}} & loc_sram_buff_w8[124][3:0]) | ({4{loc_sram_buff_w9[124][4]}} & loc_sram_buff_w9[124][3:0]) | ({4{loc_sram_buff_w10[124][4]}} & loc_sram_buff_w10[124][3:0]) | ({4{loc_sram_buff_w11[124][4]}} & loc_sram_buff_w11[124][3:0]) | ({4{loc_sram_buff_w12[124][4]}} & loc_sram_buff_w12[124][3:0]) | ({4{loc_sram_buff_w13[124][4]}} & loc_sram_buff_w13[124][3:0]) | ({4{loc_sram_buff_w14[124][4]}} & loc_sram_buff_w14[124][3:0]) | ({4{loc_sram_buff_w15[124][4]}} & loc_sram_buff_w15[124][3:0]);
	loc_rdata_buff[ 523: 520] = ({4{loc_sram_buff_w0[125][4]}} & loc_sram_buff_w0[125][3:0]) | ({4{loc_sram_buff_w1[125][4]}} & loc_sram_buff_w1[125][3:0]) | ({4{loc_sram_buff_w2[125][4]}} & loc_sram_buff_w2[125][3:0]) | ({4{loc_sram_buff_w3[125][4]}} & loc_sram_buff_w3[125][3:0]) | ({4{loc_sram_buff_w4[125][4]}} & loc_sram_buff_w4[125][3:0]) | ({4{loc_sram_buff_w5[125][4]}} & loc_sram_buff_w5[125][3:0]) | ({4{loc_sram_buff_w6[125][4]}} & loc_sram_buff_w6[125][3:0]) | ({4{loc_sram_buff_w7[125][4]}} & loc_sram_buff_w7[125][3:0]) | ({4{loc_sram_buff_w8[125][4]}} & loc_sram_buff_w8[125][3:0]) | ({4{loc_sram_buff_w9[125][4]}} & loc_sram_buff_w9[125][3:0]) | ({4{loc_sram_buff_w10[125][4]}} & loc_sram_buff_w10[125][3:0]) | ({4{loc_sram_buff_w11[125][4]}} & loc_sram_buff_w11[125][3:0]) | ({4{loc_sram_buff_w12[125][4]}} & loc_sram_buff_w12[125][3:0]) | ({4{loc_sram_buff_w13[125][4]}} & loc_sram_buff_w13[125][3:0]) | ({4{loc_sram_buff_w14[125][4]}} & loc_sram_buff_w14[125][3:0]) | ({4{loc_sram_buff_w15[125][4]}} & loc_sram_buff_w15[125][3:0]);
	loc_rdata_buff[ 519: 516] = ({4{loc_sram_buff_w0[126][4]}} & loc_sram_buff_w0[126][3:0]) | ({4{loc_sram_buff_w1[126][4]}} & loc_sram_buff_w1[126][3:0]) | ({4{loc_sram_buff_w2[126][4]}} & loc_sram_buff_w2[126][3:0]) | ({4{loc_sram_buff_w3[126][4]}} & loc_sram_buff_w3[126][3:0]) | ({4{loc_sram_buff_w4[126][4]}} & loc_sram_buff_w4[126][3:0]) | ({4{loc_sram_buff_w5[126][4]}} & loc_sram_buff_w5[126][3:0]) | ({4{loc_sram_buff_w6[126][4]}} & loc_sram_buff_w6[126][3:0]) | ({4{loc_sram_buff_w7[126][4]}} & loc_sram_buff_w7[126][3:0]) | ({4{loc_sram_buff_w8[126][4]}} & loc_sram_buff_w8[126][3:0]) | ({4{loc_sram_buff_w9[126][4]}} & loc_sram_buff_w9[126][3:0]) | ({4{loc_sram_buff_w10[126][4]}} & loc_sram_buff_w10[126][3:0]) | ({4{loc_sram_buff_w11[126][4]}} & loc_sram_buff_w11[126][3:0]) | ({4{loc_sram_buff_w12[126][4]}} & loc_sram_buff_w12[126][3:0]) | ({4{loc_sram_buff_w13[126][4]}} & loc_sram_buff_w13[126][3:0]) | ({4{loc_sram_buff_w14[126][4]}} & loc_sram_buff_w14[126][3:0]) | ({4{loc_sram_buff_w15[126][4]}} & loc_sram_buff_w15[126][3:0]);
	loc_rdata_buff[ 515: 512] = ({4{loc_sram_buff_w0[127][4]}} & loc_sram_buff_w0[127][3:0]) | ({4{loc_sram_buff_w1[127][4]}} & loc_sram_buff_w1[127][3:0]) | ({4{loc_sram_buff_w2[127][4]}} & loc_sram_buff_w2[127][3:0]) | ({4{loc_sram_buff_w3[127][4]}} & loc_sram_buff_w3[127][3:0]) | ({4{loc_sram_buff_w4[127][4]}} & loc_sram_buff_w4[127][3:0]) | ({4{loc_sram_buff_w5[127][4]}} & loc_sram_buff_w5[127][3:0]) | ({4{loc_sram_buff_w6[127][4]}} & loc_sram_buff_w6[127][3:0]) | ({4{loc_sram_buff_w7[127][4]}} & loc_sram_buff_w7[127][3:0]) | ({4{loc_sram_buff_w8[127][4]}} & loc_sram_buff_w8[127][3:0]) | ({4{loc_sram_buff_w9[127][4]}} & loc_sram_buff_w9[127][3:0]) | ({4{loc_sram_buff_w10[127][4]}} & loc_sram_buff_w10[127][3:0]) | ({4{loc_sram_buff_w11[127][4]}} & loc_sram_buff_w11[127][3:0]) | ({4{loc_sram_buff_w12[127][4]}} & loc_sram_buff_w12[127][3:0]) | ({4{loc_sram_buff_w13[127][4]}} & loc_sram_buff_w13[127][3:0]) | ({4{loc_sram_buff_w14[127][4]}} & loc_sram_buff_w14[127][3:0]) | ({4{loc_sram_buff_w15[127][4]}} & loc_sram_buff_w15[127][3:0]);
	loc_rdata_buff[ 511: 508] = ({4{loc_sram_buff_w0[128][4]}} & loc_sram_buff_w0[128][3:0]) | ({4{loc_sram_buff_w1[128][4]}} & loc_sram_buff_w1[128][3:0]) | ({4{loc_sram_buff_w2[128][4]}} & loc_sram_buff_w2[128][3:0]) | ({4{loc_sram_buff_w3[128][4]}} & loc_sram_buff_w3[128][3:0]) | ({4{loc_sram_buff_w4[128][4]}} & loc_sram_buff_w4[128][3:0]) | ({4{loc_sram_buff_w5[128][4]}} & loc_sram_buff_w5[128][3:0]) | ({4{loc_sram_buff_w6[128][4]}} & loc_sram_buff_w6[128][3:0]) | ({4{loc_sram_buff_w7[128][4]}} & loc_sram_buff_w7[128][3:0]) | ({4{loc_sram_buff_w8[128][4]}} & loc_sram_buff_w8[128][3:0]) | ({4{loc_sram_buff_w9[128][4]}} & loc_sram_buff_w9[128][3:0]) | ({4{loc_sram_buff_w10[128][4]}} & loc_sram_buff_w10[128][3:0]) | ({4{loc_sram_buff_w11[128][4]}} & loc_sram_buff_w11[128][3:0]) | ({4{loc_sram_buff_w12[128][4]}} & loc_sram_buff_w12[128][3:0]) | ({4{loc_sram_buff_w13[128][4]}} & loc_sram_buff_w13[128][3:0]) | ({4{loc_sram_buff_w14[128][4]}} & loc_sram_buff_w14[128][3:0]) | ({4{loc_sram_buff_w15[128][4]}} & loc_sram_buff_w15[128][3:0]);
	loc_rdata_buff[ 507: 504] = ({4{loc_sram_buff_w0[129][4]}} & loc_sram_buff_w0[129][3:0]) | ({4{loc_sram_buff_w1[129][4]}} & loc_sram_buff_w1[129][3:0]) | ({4{loc_sram_buff_w2[129][4]}} & loc_sram_buff_w2[129][3:0]) | ({4{loc_sram_buff_w3[129][4]}} & loc_sram_buff_w3[129][3:0]) | ({4{loc_sram_buff_w4[129][4]}} & loc_sram_buff_w4[129][3:0]) | ({4{loc_sram_buff_w5[129][4]}} & loc_sram_buff_w5[129][3:0]) | ({4{loc_sram_buff_w6[129][4]}} & loc_sram_buff_w6[129][3:0]) | ({4{loc_sram_buff_w7[129][4]}} & loc_sram_buff_w7[129][3:0]) | ({4{loc_sram_buff_w8[129][4]}} & loc_sram_buff_w8[129][3:0]) | ({4{loc_sram_buff_w9[129][4]}} & loc_sram_buff_w9[129][3:0]) | ({4{loc_sram_buff_w10[129][4]}} & loc_sram_buff_w10[129][3:0]) | ({4{loc_sram_buff_w11[129][4]}} & loc_sram_buff_w11[129][3:0]) | ({4{loc_sram_buff_w12[129][4]}} & loc_sram_buff_w12[129][3:0]) | ({4{loc_sram_buff_w13[129][4]}} & loc_sram_buff_w13[129][3:0]) | ({4{loc_sram_buff_w14[129][4]}} & loc_sram_buff_w14[129][3:0]) | ({4{loc_sram_buff_w15[129][4]}} & loc_sram_buff_w15[129][3:0]);
	loc_rdata_buff[ 503: 500] = ({4{loc_sram_buff_w0[130][4]}} & loc_sram_buff_w0[130][3:0]) | ({4{loc_sram_buff_w1[130][4]}} & loc_sram_buff_w1[130][3:0]) | ({4{loc_sram_buff_w2[130][4]}} & loc_sram_buff_w2[130][3:0]) | ({4{loc_sram_buff_w3[130][4]}} & loc_sram_buff_w3[130][3:0]) | ({4{loc_sram_buff_w4[130][4]}} & loc_sram_buff_w4[130][3:0]) | ({4{loc_sram_buff_w5[130][4]}} & loc_sram_buff_w5[130][3:0]) | ({4{loc_sram_buff_w6[130][4]}} & loc_sram_buff_w6[130][3:0]) | ({4{loc_sram_buff_w7[130][4]}} & loc_sram_buff_w7[130][3:0]) | ({4{loc_sram_buff_w8[130][4]}} & loc_sram_buff_w8[130][3:0]) | ({4{loc_sram_buff_w9[130][4]}} & loc_sram_buff_w9[130][3:0]) | ({4{loc_sram_buff_w10[130][4]}} & loc_sram_buff_w10[130][3:0]) | ({4{loc_sram_buff_w11[130][4]}} & loc_sram_buff_w11[130][3:0]) | ({4{loc_sram_buff_w12[130][4]}} & loc_sram_buff_w12[130][3:0]) | ({4{loc_sram_buff_w13[130][4]}} & loc_sram_buff_w13[130][3:0]) | ({4{loc_sram_buff_w14[130][4]}} & loc_sram_buff_w14[130][3:0]) | ({4{loc_sram_buff_w15[130][4]}} & loc_sram_buff_w15[130][3:0]);
	loc_rdata_buff[ 499: 496] = ({4{loc_sram_buff_w0[131][4]}} & loc_sram_buff_w0[131][3:0]) | ({4{loc_sram_buff_w1[131][4]}} & loc_sram_buff_w1[131][3:0]) | ({4{loc_sram_buff_w2[131][4]}} & loc_sram_buff_w2[131][3:0]) | ({4{loc_sram_buff_w3[131][4]}} & loc_sram_buff_w3[131][3:0]) | ({4{loc_sram_buff_w4[131][4]}} & loc_sram_buff_w4[131][3:0]) | ({4{loc_sram_buff_w5[131][4]}} & loc_sram_buff_w5[131][3:0]) | ({4{loc_sram_buff_w6[131][4]}} & loc_sram_buff_w6[131][3:0]) | ({4{loc_sram_buff_w7[131][4]}} & loc_sram_buff_w7[131][3:0]) | ({4{loc_sram_buff_w8[131][4]}} & loc_sram_buff_w8[131][3:0]) | ({4{loc_sram_buff_w9[131][4]}} & loc_sram_buff_w9[131][3:0]) | ({4{loc_sram_buff_w10[131][4]}} & loc_sram_buff_w10[131][3:0]) | ({4{loc_sram_buff_w11[131][4]}} & loc_sram_buff_w11[131][3:0]) | ({4{loc_sram_buff_w12[131][4]}} & loc_sram_buff_w12[131][3:0]) | ({4{loc_sram_buff_w13[131][4]}} & loc_sram_buff_w13[131][3:0]) | ({4{loc_sram_buff_w14[131][4]}} & loc_sram_buff_w14[131][3:0]) | ({4{loc_sram_buff_w15[131][4]}} & loc_sram_buff_w15[131][3:0]);
	loc_rdata_buff[ 495: 492] = ({4{loc_sram_buff_w0[132][4]}} & loc_sram_buff_w0[132][3:0]) | ({4{loc_sram_buff_w1[132][4]}} & loc_sram_buff_w1[132][3:0]) | ({4{loc_sram_buff_w2[132][4]}} & loc_sram_buff_w2[132][3:0]) | ({4{loc_sram_buff_w3[132][4]}} & loc_sram_buff_w3[132][3:0]) | ({4{loc_sram_buff_w4[132][4]}} & loc_sram_buff_w4[132][3:0]) | ({4{loc_sram_buff_w5[132][4]}} & loc_sram_buff_w5[132][3:0]) | ({4{loc_sram_buff_w6[132][4]}} & loc_sram_buff_w6[132][3:0]) | ({4{loc_sram_buff_w7[132][4]}} & loc_sram_buff_w7[132][3:0]) | ({4{loc_sram_buff_w8[132][4]}} & loc_sram_buff_w8[132][3:0]) | ({4{loc_sram_buff_w9[132][4]}} & loc_sram_buff_w9[132][3:0]) | ({4{loc_sram_buff_w10[132][4]}} & loc_sram_buff_w10[132][3:0]) | ({4{loc_sram_buff_w11[132][4]}} & loc_sram_buff_w11[132][3:0]) | ({4{loc_sram_buff_w12[132][4]}} & loc_sram_buff_w12[132][3:0]) | ({4{loc_sram_buff_w13[132][4]}} & loc_sram_buff_w13[132][3:0]) | ({4{loc_sram_buff_w14[132][4]}} & loc_sram_buff_w14[132][3:0]) | ({4{loc_sram_buff_w15[132][4]}} & loc_sram_buff_w15[132][3:0]);
	loc_rdata_buff[ 491: 488] = ({4{loc_sram_buff_w0[133][4]}} & loc_sram_buff_w0[133][3:0]) | ({4{loc_sram_buff_w1[133][4]}} & loc_sram_buff_w1[133][3:0]) | ({4{loc_sram_buff_w2[133][4]}} & loc_sram_buff_w2[133][3:0]) | ({4{loc_sram_buff_w3[133][4]}} & loc_sram_buff_w3[133][3:0]) | ({4{loc_sram_buff_w4[133][4]}} & loc_sram_buff_w4[133][3:0]) | ({4{loc_sram_buff_w5[133][4]}} & loc_sram_buff_w5[133][3:0]) | ({4{loc_sram_buff_w6[133][4]}} & loc_sram_buff_w6[133][3:0]) | ({4{loc_sram_buff_w7[133][4]}} & loc_sram_buff_w7[133][3:0]) | ({4{loc_sram_buff_w8[133][4]}} & loc_sram_buff_w8[133][3:0]) | ({4{loc_sram_buff_w9[133][4]}} & loc_sram_buff_w9[133][3:0]) | ({4{loc_sram_buff_w10[133][4]}} & loc_sram_buff_w10[133][3:0]) | ({4{loc_sram_buff_w11[133][4]}} & loc_sram_buff_w11[133][3:0]) | ({4{loc_sram_buff_w12[133][4]}} & loc_sram_buff_w12[133][3:0]) | ({4{loc_sram_buff_w13[133][4]}} & loc_sram_buff_w13[133][3:0]) | ({4{loc_sram_buff_w14[133][4]}} & loc_sram_buff_w14[133][3:0]) | ({4{loc_sram_buff_w15[133][4]}} & loc_sram_buff_w15[133][3:0]);
	loc_rdata_buff[ 487: 484] = ({4{loc_sram_buff_w0[134][4]}} & loc_sram_buff_w0[134][3:0]) | ({4{loc_sram_buff_w1[134][4]}} & loc_sram_buff_w1[134][3:0]) | ({4{loc_sram_buff_w2[134][4]}} & loc_sram_buff_w2[134][3:0]) | ({4{loc_sram_buff_w3[134][4]}} & loc_sram_buff_w3[134][3:0]) | ({4{loc_sram_buff_w4[134][4]}} & loc_sram_buff_w4[134][3:0]) | ({4{loc_sram_buff_w5[134][4]}} & loc_sram_buff_w5[134][3:0]) | ({4{loc_sram_buff_w6[134][4]}} & loc_sram_buff_w6[134][3:0]) | ({4{loc_sram_buff_w7[134][4]}} & loc_sram_buff_w7[134][3:0]) | ({4{loc_sram_buff_w8[134][4]}} & loc_sram_buff_w8[134][3:0]) | ({4{loc_sram_buff_w9[134][4]}} & loc_sram_buff_w9[134][3:0]) | ({4{loc_sram_buff_w10[134][4]}} & loc_sram_buff_w10[134][3:0]) | ({4{loc_sram_buff_w11[134][4]}} & loc_sram_buff_w11[134][3:0]) | ({4{loc_sram_buff_w12[134][4]}} & loc_sram_buff_w12[134][3:0]) | ({4{loc_sram_buff_w13[134][4]}} & loc_sram_buff_w13[134][3:0]) | ({4{loc_sram_buff_w14[134][4]}} & loc_sram_buff_w14[134][3:0]) | ({4{loc_sram_buff_w15[134][4]}} & loc_sram_buff_w15[134][3:0]);
	loc_rdata_buff[ 483: 480] = ({4{loc_sram_buff_w0[135][4]}} & loc_sram_buff_w0[135][3:0]) | ({4{loc_sram_buff_w1[135][4]}} & loc_sram_buff_w1[135][3:0]) | ({4{loc_sram_buff_w2[135][4]}} & loc_sram_buff_w2[135][3:0]) | ({4{loc_sram_buff_w3[135][4]}} & loc_sram_buff_w3[135][3:0]) | ({4{loc_sram_buff_w4[135][4]}} & loc_sram_buff_w4[135][3:0]) | ({4{loc_sram_buff_w5[135][4]}} & loc_sram_buff_w5[135][3:0]) | ({4{loc_sram_buff_w6[135][4]}} & loc_sram_buff_w6[135][3:0]) | ({4{loc_sram_buff_w7[135][4]}} & loc_sram_buff_w7[135][3:0]) | ({4{loc_sram_buff_w8[135][4]}} & loc_sram_buff_w8[135][3:0]) | ({4{loc_sram_buff_w9[135][4]}} & loc_sram_buff_w9[135][3:0]) | ({4{loc_sram_buff_w10[135][4]}} & loc_sram_buff_w10[135][3:0]) | ({4{loc_sram_buff_w11[135][4]}} & loc_sram_buff_w11[135][3:0]) | ({4{loc_sram_buff_w12[135][4]}} & loc_sram_buff_w12[135][3:0]) | ({4{loc_sram_buff_w13[135][4]}} & loc_sram_buff_w13[135][3:0]) | ({4{loc_sram_buff_w14[135][4]}} & loc_sram_buff_w14[135][3:0]) | ({4{loc_sram_buff_w15[135][4]}} & loc_sram_buff_w15[135][3:0]);
	loc_rdata_buff[ 479: 476] = ({4{loc_sram_buff_w0[136][4]}} & loc_sram_buff_w0[136][3:0]) | ({4{loc_sram_buff_w1[136][4]}} & loc_sram_buff_w1[136][3:0]) | ({4{loc_sram_buff_w2[136][4]}} & loc_sram_buff_w2[136][3:0]) | ({4{loc_sram_buff_w3[136][4]}} & loc_sram_buff_w3[136][3:0]) | ({4{loc_sram_buff_w4[136][4]}} & loc_sram_buff_w4[136][3:0]) | ({4{loc_sram_buff_w5[136][4]}} & loc_sram_buff_w5[136][3:0]) | ({4{loc_sram_buff_w6[136][4]}} & loc_sram_buff_w6[136][3:0]) | ({4{loc_sram_buff_w7[136][4]}} & loc_sram_buff_w7[136][3:0]) | ({4{loc_sram_buff_w8[136][4]}} & loc_sram_buff_w8[136][3:0]) | ({4{loc_sram_buff_w9[136][4]}} & loc_sram_buff_w9[136][3:0]) | ({4{loc_sram_buff_w10[136][4]}} & loc_sram_buff_w10[136][3:0]) | ({4{loc_sram_buff_w11[136][4]}} & loc_sram_buff_w11[136][3:0]) | ({4{loc_sram_buff_w12[136][4]}} & loc_sram_buff_w12[136][3:0]) | ({4{loc_sram_buff_w13[136][4]}} & loc_sram_buff_w13[136][3:0]) | ({4{loc_sram_buff_w14[136][4]}} & loc_sram_buff_w14[136][3:0]) | ({4{loc_sram_buff_w15[136][4]}} & loc_sram_buff_w15[136][3:0]);
	loc_rdata_buff[ 475: 472] = ({4{loc_sram_buff_w0[137][4]}} & loc_sram_buff_w0[137][3:0]) | ({4{loc_sram_buff_w1[137][4]}} & loc_sram_buff_w1[137][3:0]) | ({4{loc_sram_buff_w2[137][4]}} & loc_sram_buff_w2[137][3:0]) | ({4{loc_sram_buff_w3[137][4]}} & loc_sram_buff_w3[137][3:0]) | ({4{loc_sram_buff_w4[137][4]}} & loc_sram_buff_w4[137][3:0]) | ({4{loc_sram_buff_w5[137][4]}} & loc_sram_buff_w5[137][3:0]) | ({4{loc_sram_buff_w6[137][4]}} & loc_sram_buff_w6[137][3:0]) | ({4{loc_sram_buff_w7[137][4]}} & loc_sram_buff_w7[137][3:0]) | ({4{loc_sram_buff_w8[137][4]}} & loc_sram_buff_w8[137][3:0]) | ({4{loc_sram_buff_w9[137][4]}} & loc_sram_buff_w9[137][3:0]) | ({4{loc_sram_buff_w10[137][4]}} & loc_sram_buff_w10[137][3:0]) | ({4{loc_sram_buff_w11[137][4]}} & loc_sram_buff_w11[137][3:0]) | ({4{loc_sram_buff_w12[137][4]}} & loc_sram_buff_w12[137][3:0]) | ({4{loc_sram_buff_w13[137][4]}} & loc_sram_buff_w13[137][3:0]) | ({4{loc_sram_buff_w14[137][4]}} & loc_sram_buff_w14[137][3:0]) | ({4{loc_sram_buff_w15[137][4]}} & loc_sram_buff_w15[137][3:0]);
	loc_rdata_buff[ 471: 468] = ({4{loc_sram_buff_w0[138][4]}} & loc_sram_buff_w0[138][3:0]) | ({4{loc_sram_buff_w1[138][4]}} & loc_sram_buff_w1[138][3:0]) | ({4{loc_sram_buff_w2[138][4]}} & loc_sram_buff_w2[138][3:0]) | ({4{loc_sram_buff_w3[138][4]}} & loc_sram_buff_w3[138][3:0]) | ({4{loc_sram_buff_w4[138][4]}} & loc_sram_buff_w4[138][3:0]) | ({4{loc_sram_buff_w5[138][4]}} & loc_sram_buff_w5[138][3:0]) | ({4{loc_sram_buff_w6[138][4]}} & loc_sram_buff_w6[138][3:0]) | ({4{loc_sram_buff_w7[138][4]}} & loc_sram_buff_w7[138][3:0]) | ({4{loc_sram_buff_w8[138][4]}} & loc_sram_buff_w8[138][3:0]) | ({4{loc_sram_buff_w9[138][4]}} & loc_sram_buff_w9[138][3:0]) | ({4{loc_sram_buff_w10[138][4]}} & loc_sram_buff_w10[138][3:0]) | ({4{loc_sram_buff_w11[138][4]}} & loc_sram_buff_w11[138][3:0]) | ({4{loc_sram_buff_w12[138][4]}} & loc_sram_buff_w12[138][3:0]) | ({4{loc_sram_buff_w13[138][4]}} & loc_sram_buff_w13[138][3:0]) | ({4{loc_sram_buff_w14[138][4]}} & loc_sram_buff_w14[138][3:0]) | ({4{loc_sram_buff_w15[138][4]}} & loc_sram_buff_w15[138][3:0]);
	loc_rdata_buff[ 467: 464] = ({4{loc_sram_buff_w0[139][4]}} & loc_sram_buff_w0[139][3:0]) | ({4{loc_sram_buff_w1[139][4]}} & loc_sram_buff_w1[139][3:0]) | ({4{loc_sram_buff_w2[139][4]}} & loc_sram_buff_w2[139][3:0]) | ({4{loc_sram_buff_w3[139][4]}} & loc_sram_buff_w3[139][3:0]) | ({4{loc_sram_buff_w4[139][4]}} & loc_sram_buff_w4[139][3:0]) | ({4{loc_sram_buff_w5[139][4]}} & loc_sram_buff_w5[139][3:0]) | ({4{loc_sram_buff_w6[139][4]}} & loc_sram_buff_w6[139][3:0]) | ({4{loc_sram_buff_w7[139][4]}} & loc_sram_buff_w7[139][3:0]) | ({4{loc_sram_buff_w8[139][4]}} & loc_sram_buff_w8[139][3:0]) | ({4{loc_sram_buff_w9[139][4]}} & loc_sram_buff_w9[139][3:0]) | ({4{loc_sram_buff_w10[139][4]}} & loc_sram_buff_w10[139][3:0]) | ({4{loc_sram_buff_w11[139][4]}} & loc_sram_buff_w11[139][3:0]) | ({4{loc_sram_buff_w12[139][4]}} & loc_sram_buff_w12[139][3:0]) | ({4{loc_sram_buff_w13[139][4]}} & loc_sram_buff_w13[139][3:0]) | ({4{loc_sram_buff_w14[139][4]}} & loc_sram_buff_w14[139][3:0]) | ({4{loc_sram_buff_w15[139][4]}} & loc_sram_buff_w15[139][3:0]);
	loc_rdata_buff[ 463: 460] = ({4{loc_sram_buff_w0[140][4]}} & loc_sram_buff_w0[140][3:0]) | ({4{loc_sram_buff_w1[140][4]}} & loc_sram_buff_w1[140][3:0]) | ({4{loc_sram_buff_w2[140][4]}} & loc_sram_buff_w2[140][3:0]) | ({4{loc_sram_buff_w3[140][4]}} & loc_sram_buff_w3[140][3:0]) | ({4{loc_sram_buff_w4[140][4]}} & loc_sram_buff_w4[140][3:0]) | ({4{loc_sram_buff_w5[140][4]}} & loc_sram_buff_w5[140][3:0]) | ({4{loc_sram_buff_w6[140][4]}} & loc_sram_buff_w6[140][3:0]) | ({4{loc_sram_buff_w7[140][4]}} & loc_sram_buff_w7[140][3:0]) | ({4{loc_sram_buff_w8[140][4]}} & loc_sram_buff_w8[140][3:0]) | ({4{loc_sram_buff_w9[140][4]}} & loc_sram_buff_w9[140][3:0]) | ({4{loc_sram_buff_w10[140][4]}} & loc_sram_buff_w10[140][3:0]) | ({4{loc_sram_buff_w11[140][4]}} & loc_sram_buff_w11[140][3:0]) | ({4{loc_sram_buff_w12[140][4]}} & loc_sram_buff_w12[140][3:0]) | ({4{loc_sram_buff_w13[140][4]}} & loc_sram_buff_w13[140][3:0]) | ({4{loc_sram_buff_w14[140][4]}} & loc_sram_buff_w14[140][3:0]) | ({4{loc_sram_buff_w15[140][4]}} & loc_sram_buff_w15[140][3:0]);
	loc_rdata_buff[ 459: 456] = ({4{loc_sram_buff_w0[141][4]}} & loc_sram_buff_w0[141][3:0]) | ({4{loc_sram_buff_w1[141][4]}} & loc_sram_buff_w1[141][3:0]) | ({4{loc_sram_buff_w2[141][4]}} & loc_sram_buff_w2[141][3:0]) | ({4{loc_sram_buff_w3[141][4]}} & loc_sram_buff_w3[141][3:0]) | ({4{loc_sram_buff_w4[141][4]}} & loc_sram_buff_w4[141][3:0]) | ({4{loc_sram_buff_w5[141][4]}} & loc_sram_buff_w5[141][3:0]) | ({4{loc_sram_buff_w6[141][4]}} & loc_sram_buff_w6[141][3:0]) | ({4{loc_sram_buff_w7[141][4]}} & loc_sram_buff_w7[141][3:0]) | ({4{loc_sram_buff_w8[141][4]}} & loc_sram_buff_w8[141][3:0]) | ({4{loc_sram_buff_w9[141][4]}} & loc_sram_buff_w9[141][3:0]) | ({4{loc_sram_buff_w10[141][4]}} & loc_sram_buff_w10[141][3:0]) | ({4{loc_sram_buff_w11[141][4]}} & loc_sram_buff_w11[141][3:0]) | ({4{loc_sram_buff_w12[141][4]}} & loc_sram_buff_w12[141][3:0]) | ({4{loc_sram_buff_w13[141][4]}} & loc_sram_buff_w13[141][3:0]) | ({4{loc_sram_buff_w14[141][4]}} & loc_sram_buff_w14[141][3:0]) | ({4{loc_sram_buff_w15[141][4]}} & loc_sram_buff_w15[141][3:0]);
	loc_rdata_buff[ 455: 452] = ({4{loc_sram_buff_w0[142][4]}} & loc_sram_buff_w0[142][3:0]) | ({4{loc_sram_buff_w1[142][4]}} & loc_sram_buff_w1[142][3:0]) | ({4{loc_sram_buff_w2[142][4]}} & loc_sram_buff_w2[142][3:0]) | ({4{loc_sram_buff_w3[142][4]}} & loc_sram_buff_w3[142][3:0]) | ({4{loc_sram_buff_w4[142][4]}} & loc_sram_buff_w4[142][3:0]) | ({4{loc_sram_buff_w5[142][4]}} & loc_sram_buff_w5[142][3:0]) | ({4{loc_sram_buff_w6[142][4]}} & loc_sram_buff_w6[142][3:0]) | ({4{loc_sram_buff_w7[142][4]}} & loc_sram_buff_w7[142][3:0]) | ({4{loc_sram_buff_w8[142][4]}} & loc_sram_buff_w8[142][3:0]) | ({4{loc_sram_buff_w9[142][4]}} & loc_sram_buff_w9[142][3:0]) | ({4{loc_sram_buff_w10[142][4]}} & loc_sram_buff_w10[142][3:0]) | ({4{loc_sram_buff_w11[142][4]}} & loc_sram_buff_w11[142][3:0]) | ({4{loc_sram_buff_w12[142][4]}} & loc_sram_buff_w12[142][3:0]) | ({4{loc_sram_buff_w13[142][4]}} & loc_sram_buff_w13[142][3:0]) | ({4{loc_sram_buff_w14[142][4]}} & loc_sram_buff_w14[142][3:0]) | ({4{loc_sram_buff_w15[142][4]}} & loc_sram_buff_w15[142][3:0]);
	loc_rdata_buff[ 451: 448] = ({4{loc_sram_buff_w0[143][4]}} & loc_sram_buff_w0[143][3:0]) | ({4{loc_sram_buff_w1[143][4]}} & loc_sram_buff_w1[143][3:0]) | ({4{loc_sram_buff_w2[143][4]}} & loc_sram_buff_w2[143][3:0]) | ({4{loc_sram_buff_w3[143][4]}} & loc_sram_buff_w3[143][3:0]) | ({4{loc_sram_buff_w4[143][4]}} & loc_sram_buff_w4[143][3:0]) | ({4{loc_sram_buff_w5[143][4]}} & loc_sram_buff_w5[143][3:0]) | ({4{loc_sram_buff_w6[143][4]}} & loc_sram_buff_w6[143][3:0]) | ({4{loc_sram_buff_w7[143][4]}} & loc_sram_buff_w7[143][3:0]) | ({4{loc_sram_buff_w8[143][4]}} & loc_sram_buff_w8[143][3:0]) | ({4{loc_sram_buff_w9[143][4]}} & loc_sram_buff_w9[143][3:0]) | ({4{loc_sram_buff_w10[143][4]}} & loc_sram_buff_w10[143][3:0]) | ({4{loc_sram_buff_w11[143][4]}} & loc_sram_buff_w11[143][3:0]) | ({4{loc_sram_buff_w12[143][4]}} & loc_sram_buff_w12[143][3:0]) | ({4{loc_sram_buff_w13[143][4]}} & loc_sram_buff_w13[143][3:0]) | ({4{loc_sram_buff_w14[143][4]}} & loc_sram_buff_w14[143][3:0]) | ({4{loc_sram_buff_w15[143][4]}} & loc_sram_buff_w15[143][3:0]);
	loc_rdata_buff[ 447: 444] = ({4{loc_sram_buff_w0[144][4]}} & loc_sram_buff_w0[144][3:0]) | ({4{loc_sram_buff_w1[144][4]}} & loc_sram_buff_w1[144][3:0]) | ({4{loc_sram_buff_w2[144][4]}} & loc_sram_buff_w2[144][3:0]) | ({4{loc_sram_buff_w3[144][4]}} & loc_sram_buff_w3[144][3:0]) | ({4{loc_sram_buff_w4[144][4]}} & loc_sram_buff_w4[144][3:0]) | ({4{loc_sram_buff_w5[144][4]}} & loc_sram_buff_w5[144][3:0]) | ({4{loc_sram_buff_w6[144][4]}} & loc_sram_buff_w6[144][3:0]) | ({4{loc_sram_buff_w7[144][4]}} & loc_sram_buff_w7[144][3:0]) | ({4{loc_sram_buff_w8[144][4]}} & loc_sram_buff_w8[144][3:0]) | ({4{loc_sram_buff_w9[144][4]}} & loc_sram_buff_w9[144][3:0]) | ({4{loc_sram_buff_w10[144][4]}} & loc_sram_buff_w10[144][3:0]) | ({4{loc_sram_buff_w11[144][4]}} & loc_sram_buff_w11[144][3:0]) | ({4{loc_sram_buff_w12[144][4]}} & loc_sram_buff_w12[144][3:0]) | ({4{loc_sram_buff_w13[144][4]}} & loc_sram_buff_w13[144][3:0]) | ({4{loc_sram_buff_w14[144][4]}} & loc_sram_buff_w14[144][3:0]) | ({4{loc_sram_buff_w15[144][4]}} & loc_sram_buff_w15[144][3:0]);
	loc_rdata_buff[ 443: 440] = ({4{loc_sram_buff_w0[145][4]}} & loc_sram_buff_w0[145][3:0]) | ({4{loc_sram_buff_w1[145][4]}} & loc_sram_buff_w1[145][3:0]) | ({4{loc_sram_buff_w2[145][4]}} & loc_sram_buff_w2[145][3:0]) | ({4{loc_sram_buff_w3[145][4]}} & loc_sram_buff_w3[145][3:0]) | ({4{loc_sram_buff_w4[145][4]}} & loc_sram_buff_w4[145][3:0]) | ({4{loc_sram_buff_w5[145][4]}} & loc_sram_buff_w5[145][3:0]) | ({4{loc_sram_buff_w6[145][4]}} & loc_sram_buff_w6[145][3:0]) | ({4{loc_sram_buff_w7[145][4]}} & loc_sram_buff_w7[145][3:0]) | ({4{loc_sram_buff_w8[145][4]}} & loc_sram_buff_w8[145][3:0]) | ({4{loc_sram_buff_w9[145][4]}} & loc_sram_buff_w9[145][3:0]) | ({4{loc_sram_buff_w10[145][4]}} & loc_sram_buff_w10[145][3:0]) | ({4{loc_sram_buff_w11[145][4]}} & loc_sram_buff_w11[145][3:0]) | ({4{loc_sram_buff_w12[145][4]}} & loc_sram_buff_w12[145][3:0]) | ({4{loc_sram_buff_w13[145][4]}} & loc_sram_buff_w13[145][3:0]) | ({4{loc_sram_buff_w14[145][4]}} & loc_sram_buff_w14[145][3:0]) | ({4{loc_sram_buff_w15[145][4]}} & loc_sram_buff_w15[145][3:0]);
	loc_rdata_buff[ 439: 436] = ({4{loc_sram_buff_w0[146][4]}} & loc_sram_buff_w0[146][3:0]) | ({4{loc_sram_buff_w1[146][4]}} & loc_sram_buff_w1[146][3:0]) | ({4{loc_sram_buff_w2[146][4]}} & loc_sram_buff_w2[146][3:0]) | ({4{loc_sram_buff_w3[146][4]}} & loc_sram_buff_w3[146][3:0]) | ({4{loc_sram_buff_w4[146][4]}} & loc_sram_buff_w4[146][3:0]) | ({4{loc_sram_buff_w5[146][4]}} & loc_sram_buff_w5[146][3:0]) | ({4{loc_sram_buff_w6[146][4]}} & loc_sram_buff_w6[146][3:0]) | ({4{loc_sram_buff_w7[146][4]}} & loc_sram_buff_w7[146][3:0]) | ({4{loc_sram_buff_w8[146][4]}} & loc_sram_buff_w8[146][3:0]) | ({4{loc_sram_buff_w9[146][4]}} & loc_sram_buff_w9[146][3:0]) | ({4{loc_sram_buff_w10[146][4]}} & loc_sram_buff_w10[146][3:0]) | ({4{loc_sram_buff_w11[146][4]}} & loc_sram_buff_w11[146][3:0]) | ({4{loc_sram_buff_w12[146][4]}} & loc_sram_buff_w12[146][3:0]) | ({4{loc_sram_buff_w13[146][4]}} & loc_sram_buff_w13[146][3:0]) | ({4{loc_sram_buff_w14[146][4]}} & loc_sram_buff_w14[146][3:0]) | ({4{loc_sram_buff_w15[146][4]}} & loc_sram_buff_w15[146][3:0]);
	loc_rdata_buff[ 435: 432] = ({4{loc_sram_buff_w0[147][4]}} & loc_sram_buff_w0[147][3:0]) | ({4{loc_sram_buff_w1[147][4]}} & loc_sram_buff_w1[147][3:0]) | ({4{loc_sram_buff_w2[147][4]}} & loc_sram_buff_w2[147][3:0]) | ({4{loc_sram_buff_w3[147][4]}} & loc_sram_buff_w3[147][3:0]) | ({4{loc_sram_buff_w4[147][4]}} & loc_sram_buff_w4[147][3:0]) | ({4{loc_sram_buff_w5[147][4]}} & loc_sram_buff_w5[147][3:0]) | ({4{loc_sram_buff_w6[147][4]}} & loc_sram_buff_w6[147][3:0]) | ({4{loc_sram_buff_w7[147][4]}} & loc_sram_buff_w7[147][3:0]) | ({4{loc_sram_buff_w8[147][4]}} & loc_sram_buff_w8[147][3:0]) | ({4{loc_sram_buff_w9[147][4]}} & loc_sram_buff_w9[147][3:0]) | ({4{loc_sram_buff_w10[147][4]}} & loc_sram_buff_w10[147][3:0]) | ({4{loc_sram_buff_w11[147][4]}} & loc_sram_buff_w11[147][3:0]) | ({4{loc_sram_buff_w12[147][4]}} & loc_sram_buff_w12[147][3:0]) | ({4{loc_sram_buff_w13[147][4]}} & loc_sram_buff_w13[147][3:0]) | ({4{loc_sram_buff_w14[147][4]}} & loc_sram_buff_w14[147][3:0]) | ({4{loc_sram_buff_w15[147][4]}} & loc_sram_buff_w15[147][3:0]);
	loc_rdata_buff[ 431: 428] = ({4{loc_sram_buff_w0[148][4]}} & loc_sram_buff_w0[148][3:0]) | ({4{loc_sram_buff_w1[148][4]}} & loc_sram_buff_w1[148][3:0]) | ({4{loc_sram_buff_w2[148][4]}} & loc_sram_buff_w2[148][3:0]) | ({4{loc_sram_buff_w3[148][4]}} & loc_sram_buff_w3[148][3:0]) | ({4{loc_sram_buff_w4[148][4]}} & loc_sram_buff_w4[148][3:0]) | ({4{loc_sram_buff_w5[148][4]}} & loc_sram_buff_w5[148][3:0]) | ({4{loc_sram_buff_w6[148][4]}} & loc_sram_buff_w6[148][3:0]) | ({4{loc_sram_buff_w7[148][4]}} & loc_sram_buff_w7[148][3:0]) | ({4{loc_sram_buff_w8[148][4]}} & loc_sram_buff_w8[148][3:0]) | ({4{loc_sram_buff_w9[148][4]}} & loc_sram_buff_w9[148][3:0]) | ({4{loc_sram_buff_w10[148][4]}} & loc_sram_buff_w10[148][3:0]) | ({4{loc_sram_buff_w11[148][4]}} & loc_sram_buff_w11[148][3:0]) | ({4{loc_sram_buff_w12[148][4]}} & loc_sram_buff_w12[148][3:0]) | ({4{loc_sram_buff_w13[148][4]}} & loc_sram_buff_w13[148][3:0]) | ({4{loc_sram_buff_w14[148][4]}} & loc_sram_buff_w14[148][3:0]) | ({4{loc_sram_buff_w15[148][4]}} & loc_sram_buff_w15[148][3:0]);
	loc_rdata_buff[ 427: 424] = ({4{loc_sram_buff_w0[149][4]}} & loc_sram_buff_w0[149][3:0]) | ({4{loc_sram_buff_w1[149][4]}} & loc_sram_buff_w1[149][3:0]) | ({4{loc_sram_buff_w2[149][4]}} & loc_sram_buff_w2[149][3:0]) | ({4{loc_sram_buff_w3[149][4]}} & loc_sram_buff_w3[149][3:0]) | ({4{loc_sram_buff_w4[149][4]}} & loc_sram_buff_w4[149][3:0]) | ({4{loc_sram_buff_w5[149][4]}} & loc_sram_buff_w5[149][3:0]) | ({4{loc_sram_buff_w6[149][4]}} & loc_sram_buff_w6[149][3:0]) | ({4{loc_sram_buff_w7[149][4]}} & loc_sram_buff_w7[149][3:0]) | ({4{loc_sram_buff_w8[149][4]}} & loc_sram_buff_w8[149][3:0]) | ({4{loc_sram_buff_w9[149][4]}} & loc_sram_buff_w9[149][3:0]) | ({4{loc_sram_buff_w10[149][4]}} & loc_sram_buff_w10[149][3:0]) | ({4{loc_sram_buff_w11[149][4]}} & loc_sram_buff_w11[149][3:0]) | ({4{loc_sram_buff_w12[149][4]}} & loc_sram_buff_w12[149][3:0]) | ({4{loc_sram_buff_w13[149][4]}} & loc_sram_buff_w13[149][3:0]) | ({4{loc_sram_buff_w14[149][4]}} & loc_sram_buff_w14[149][3:0]) | ({4{loc_sram_buff_w15[149][4]}} & loc_sram_buff_w15[149][3:0]);
	loc_rdata_buff[ 423: 420] = ({4{loc_sram_buff_w0[150][4]}} & loc_sram_buff_w0[150][3:0]) | ({4{loc_sram_buff_w1[150][4]}} & loc_sram_buff_w1[150][3:0]) | ({4{loc_sram_buff_w2[150][4]}} & loc_sram_buff_w2[150][3:0]) | ({4{loc_sram_buff_w3[150][4]}} & loc_sram_buff_w3[150][3:0]) | ({4{loc_sram_buff_w4[150][4]}} & loc_sram_buff_w4[150][3:0]) | ({4{loc_sram_buff_w5[150][4]}} & loc_sram_buff_w5[150][3:0]) | ({4{loc_sram_buff_w6[150][4]}} & loc_sram_buff_w6[150][3:0]) | ({4{loc_sram_buff_w7[150][4]}} & loc_sram_buff_w7[150][3:0]) | ({4{loc_sram_buff_w8[150][4]}} & loc_sram_buff_w8[150][3:0]) | ({4{loc_sram_buff_w9[150][4]}} & loc_sram_buff_w9[150][3:0]) | ({4{loc_sram_buff_w10[150][4]}} & loc_sram_buff_w10[150][3:0]) | ({4{loc_sram_buff_w11[150][4]}} & loc_sram_buff_w11[150][3:0]) | ({4{loc_sram_buff_w12[150][4]}} & loc_sram_buff_w12[150][3:0]) | ({4{loc_sram_buff_w13[150][4]}} & loc_sram_buff_w13[150][3:0]) | ({4{loc_sram_buff_w14[150][4]}} & loc_sram_buff_w14[150][3:0]) | ({4{loc_sram_buff_w15[150][4]}} & loc_sram_buff_w15[150][3:0]);
	loc_rdata_buff[ 419: 416] = ({4{loc_sram_buff_w0[151][4]}} & loc_sram_buff_w0[151][3:0]) | ({4{loc_sram_buff_w1[151][4]}} & loc_sram_buff_w1[151][3:0]) | ({4{loc_sram_buff_w2[151][4]}} & loc_sram_buff_w2[151][3:0]) | ({4{loc_sram_buff_w3[151][4]}} & loc_sram_buff_w3[151][3:0]) | ({4{loc_sram_buff_w4[151][4]}} & loc_sram_buff_w4[151][3:0]) | ({4{loc_sram_buff_w5[151][4]}} & loc_sram_buff_w5[151][3:0]) | ({4{loc_sram_buff_w6[151][4]}} & loc_sram_buff_w6[151][3:0]) | ({4{loc_sram_buff_w7[151][4]}} & loc_sram_buff_w7[151][3:0]) | ({4{loc_sram_buff_w8[151][4]}} & loc_sram_buff_w8[151][3:0]) | ({4{loc_sram_buff_w9[151][4]}} & loc_sram_buff_w9[151][3:0]) | ({4{loc_sram_buff_w10[151][4]}} & loc_sram_buff_w10[151][3:0]) | ({4{loc_sram_buff_w11[151][4]}} & loc_sram_buff_w11[151][3:0]) | ({4{loc_sram_buff_w12[151][4]}} & loc_sram_buff_w12[151][3:0]) | ({4{loc_sram_buff_w13[151][4]}} & loc_sram_buff_w13[151][3:0]) | ({4{loc_sram_buff_w14[151][4]}} & loc_sram_buff_w14[151][3:0]) | ({4{loc_sram_buff_w15[151][4]}} & loc_sram_buff_w15[151][3:0]);
	loc_rdata_buff[ 415: 412] = ({4{loc_sram_buff_w0[152][4]}} & loc_sram_buff_w0[152][3:0]) | ({4{loc_sram_buff_w1[152][4]}} & loc_sram_buff_w1[152][3:0]) | ({4{loc_sram_buff_w2[152][4]}} & loc_sram_buff_w2[152][3:0]) | ({4{loc_sram_buff_w3[152][4]}} & loc_sram_buff_w3[152][3:0]) | ({4{loc_sram_buff_w4[152][4]}} & loc_sram_buff_w4[152][3:0]) | ({4{loc_sram_buff_w5[152][4]}} & loc_sram_buff_w5[152][3:0]) | ({4{loc_sram_buff_w6[152][4]}} & loc_sram_buff_w6[152][3:0]) | ({4{loc_sram_buff_w7[152][4]}} & loc_sram_buff_w7[152][3:0]) | ({4{loc_sram_buff_w8[152][4]}} & loc_sram_buff_w8[152][3:0]) | ({4{loc_sram_buff_w9[152][4]}} & loc_sram_buff_w9[152][3:0]) | ({4{loc_sram_buff_w10[152][4]}} & loc_sram_buff_w10[152][3:0]) | ({4{loc_sram_buff_w11[152][4]}} & loc_sram_buff_w11[152][3:0]) | ({4{loc_sram_buff_w12[152][4]}} & loc_sram_buff_w12[152][3:0]) | ({4{loc_sram_buff_w13[152][4]}} & loc_sram_buff_w13[152][3:0]) | ({4{loc_sram_buff_w14[152][4]}} & loc_sram_buff_w14[152][3:0]) | ({4{loc_sram_buff_w15[152][4]}} & loc_sram_buff_w15[152][3:0]);
	loc_rdata_buff[ 411: 408] = ({4{loc_sram_buff_w0[153][4]}} & loc_sram_buff_w0[153][3:0]) | ({4{loc_sram_buff_w1[153][4]}} & loc_sram_buff_w1[153][3:0]) | ({4{loc_sram_buff_w2[153][4]}} & loc_sram_buff_w2[153][3:0]) | ({4{loc_sram_buff_w3[153][4]}} & loc_sram_buff_w3[153][3:0]) | ({4{loc_sram_buff_w4[153][4]}} & loc_sram_buff_w4[153][3:0]) | ({4{loc_sram_buff_w5[153][4]}} & loc_sram_buff_w5[153][3:0]) | ({4{loc_sram_buff_w6[153][4]}} & loc_sram_buff_w6[153][3:0]) | ({4{loc_sram_buff_w7[153][4]}} & loc_sram_buff_w7[153][3:0]) | ({4{loc_sram_buff_w8[153][4]}} & loc_sram_buff_w8[153][3:0]) | ({4{loc_sram_buff_w9[153][4]}} & loc_sram_buff_w9[153][3:0]) | ({4{loc_sram_buff_w10[153][4]}} & loc_sram_buff_w10[153][3:0]) | ({4{loc_sram_buff_w11[153][4]}} & loc_sram_buff_w11[153][3:0]) | ({4{loc_sram_buff_w12[153][4]}} & loc_sram_buff_w12[153][3:0]) | ({4{loc_sram_buff_w13[153][4]}} & loc_sram_buff_w13[153][3:0]) | ({4{loc_sram_buff_w14[153][4]}} & loc_sram_buff_w14[153][3:0]) | ({4{loc_sram_buff_w15[153][4]}} & loc_sram_buff_w15[153][3:0]);
	loc_rdata_buff[ 407: 404] = ({4{loc_sram_buff_w0[154][4]}} & loc_sram_buff_w0[154][3:0]) | ({4{loc_sram_buff_w1[154][4]}} & loc_sram_buff_w1[154][3:0]) | ({4{loc_sram_buff_w2[154][4]}} & loc_sram_buff_w2[154][3:0]) | ({4{loc_sram_buff_w3[154][4]}} & loc_sram_buff_w3[154][3:0]) | ({4{loc_sram_buff_w4[154][4]}} & loc_sram_buff_w4[154][3:0]) | ({4{loc_sram_buff_w5[154][4]}} & loc_sram_buff_w5[154][3:0]) | ({4{loc_sram_buff_w6[154][4]}} & loc_sram_buff_w6[154][3:0]) | ({4{loc_sram_buff_w7[154][4]}} & loc_sram_buff_w7[154][3:0]) | ({4{loc_sram_buff_w8[154][4]}} & loc_sram_buff_w8[154][3:0]) | ({4{loc_sram_buff_w9[154][4]}} & loc_sram_buff_w9[154][3:0]) | ({4{loc_sram_buff_w10[154][4]}} & loc_sram_buff_w10[154][3:0]) | ({4{loc_sram_buff_w11[154][4]}} & loc_sram_buff_w11[154][3:0]) | ({4{loc_sram_buff_w12[154][4]}} & loc_sram_buff_w12[154][3:0]) | ({4{loc_sram_buff_w13[154][4]}} & loc_sram_buff_w13[154][3:0]) | ({4{loc_sram_buff_w14[154][4]}} & loc_sram_buff_w14[154][3:0]) | ({4{loc_sram_buff_w15[154][4]}} & loc_sram_buff_w15[154][3:0]);
	loc_rdata_buff[ 403: 400] = ({4{loc_sram_buff_w0[155][4]}} & loc_sram_buff_w0[155][3:0]) | ({4{loc_sram_buff_w1[155][4]}} & loc_sram_buff_w1[155][3:0]) | ({4{loc_sram_buff_w2[155][4]}} & loc_sram_buff_w2[155][3:0]) | ({4{loc_sram_buff_w3[155][4]}} & loc_sram_buff_w3[155][3:0]) | ({4{loc_sram_buff_w4[155][4]}} & loc_sram_buff_w4[155][3:0]) | ({4{loc_sram_buff_w5[155][4]}} & loc_sram_buff_w5[155][3:0]) | ({4{loc_sram_buff_w6[155][4]}} & loc_sram_buff_w6[155][3:0]) | ({4{loc_sram_buff_w7[155][4]}} & loc_sram_buff_w7[155][3:0]) | ({4{loc_sram_buff_w8[155][4]}} & loc_sram_buff_w8[155][3:0]) | ({4{loc_sram_buff_w9[155][4]}} & loc_sram_buff_w9[155][3:0]) | ({4{loc_sram_buff_w10[155][4]}} & loc_sram_buff_w10[155][3:0]) | ({4{loc_sram_buff_w11[155][4]}} & loc_sram_buff_w11[155][3:0]) | ({4{loc_sram_buff_w12[155][4]}} & loc_sram_buff_w12[155][3:0]) | ({4{loc_sram_buff_w13[155][4]}} & loc_sram_buff_w13[155][3:0]) | ({4{loc_sram_buff_w14[155][4]}} & loc_sram_buff_w14[155][3:0]) | ({4{loc_sram_buff_w15[155][4]}} & loc_sram_buff_w15[155][3:0]);
	loc_rdata_buff[ 399: 396] = ({4{loc_sram_buff_w0[156][4]}} & loc_sram_buff_w0[156][3:0]) | ({4{loc_sram_buff_w1[156][4]}} & loc_sram_buff_w1[156][3:0]) | ({4{loc_sram_buff_w2[156][4]}} & loc_sram_buff_w2[156][3:0]) | ({4{loc_sram_buff_w3[156][4]}} & loc_sram_buff_w3[156][3:0]) | ({4{loc_sram_buff_w4[156][4]}} & loc_sram_buff_w4[156][3:0]) | ({4{loc_sram_buff_w5[156][4]}} & loc_sram_buff_w5[156][3:0]) | ({4{loc_sram_buff_w6[156][4]}} & loc_sram_buff_w6[156][3:0]) | ({4{loc_sram_buff_w7[156][4]}} & loc_sram_buff_w7[156][3:0]) | ({4{loc_sram_buff_w8[156][4]}} & loc_sram_buff_w8[156][3:0]) | ({4{loc_sram_buff_w9[156][4]}} & loc_sram_buff_w9[156][3:0]) | ({4{loc_sram_buff_w10[156][4]}} & loc_sram_buff_w10[156][3:0]) | ({4{loc_sram_buff_w11[156][4]}} & loc_sram_buff_w11[156][3:0]) | ({4{loc_sram_buff_w12[156][4]}} & loc_sram_buff_w12[156][3:0]) | ({4{loc_sram_buff_w13[156][4]}} & loc_sram_buff_w13[156][3:0]) | ({4{loc_sram_buff_w14[156][4]}} & loc_sram_buff_w14[156][3:0]) | ({4{loc_sram_buff_w15[156][4]}} & loc_sram_buff_w15[156][3:0]);
	loc_rdata_buff[ 395: 392] = ({4{loc_sram_buff_w0[157][4]}} & loc_sram_buff_w0[157][3:0]) | ({4{loc_sram_buff_w1[157][4]}} & loc_sram_buff_w1[157][3:0]) | ({4{loc_sram_buff_w2[157][4]}} & loc_sram_buff_w2[157][3:0]) | ({4{loc_sram_buff_w3[157][4]}} & loc_sram_buff_w3[157][3:0]) | ({4{loc_sram_buff_w4[157][4]}} & loc_sram_buff_w4[157][3:0]) | ({4{loc_sram_buff_w5[157][4]}} & loc_sram_buff_w5[157][3:0]) | ({4{loc_sram_buff_w6[157][4]}} & loc_sram_buff_w6[157][3:0]) | ({4{loc_sram_buff_w7[157][4]}} & loc_sram_buff_w7[157][3:0]) | ({4{loc_sram_buff_w8[157][4]}} & loc_sram_buff_w8[157][3:0]) | ({4{loc_sram_buff_w9[157][4]}} & loc_sram_buff_w9[157][3:0]) | ({4{loc_sram_buff_w10[157][4]}} & loc_sram_buff_w10[157][3:0]) | ({4{loc_sram_buff_w11[157][4]}} & loc_sram_buff_w11[157][3:0]) | ({4{loc_sram_buff_w12[157][4]}} & loc_sram_buff_w12[157][3:0]) | ({4{loc_sram_buff_w13[157][4]}} & loc_sram_buff_w13[157][3:0]) | ({4{loc_sram_buff_w14[157][4]}} & loc_sram_buff_w14[157][3:0]) | ({4{loc_sram_buff_w15[157][4]}} & loc_sram_buff_w15[157][3:0]);
	loc_rdata_buff[ 391: 388] = ({4{loc_sram_buff_w0[158][4]}} & loc_sram_buff_w0[158][3:0]) | ({4{loc_sram_buff_w1[158][4]}} & loc_sram_buff_w1[158][3:0]) | ({4{loc_sram_buff_w2[158][4]}} & loc_sram_buff_w2[158][3:0]) | ({4{loc_sram_buff_w3[158][4]}} & loc_sram_buff_w3[158][3:0]) | ({4{loc_sram_buff_w4[158][4]}} & loc_sram_buff_w4[158][3:0]) | ({4{loc_sram_buff_w5[158][4]}} & loc_sram_buff_w5[158][3:0]) | ({4{loc_sram_buff_w6[158][4]}} & loc_sram_buff_w6[158][3:0]) | ({4{loc_sram_buff_w7[158][4]}} & loc_sram_buff_w7[158][3:0]) | ({4{loc_sram_buff_w8[158][4]}} & loc_sram_buff_w8[158][3:0]) | ({4{loc_sram_buff_w9[158][4]}} & loc_sram_buff_w9[158][3:0]) | ({4{loc_sram_buff_w10[158][4]}} & loc_sram_buff_w10[158][3:0]) | ({4{loc_sram_buff_w11[158][4]}} & loc_sram_buff_w11[158][3:0]) | ({4{loc_sram_buff_w12[158][4]}} & loc_sram_buff_w12[158][3:0]) | ({4{loc_sram_buff_w13[158][4]}} & loc_sram_buff_w13[158][3:0]) | ({4{loc_sram_buff_w14[158][4]}} & loc_sram_buff_w14[158][3:0]) | ({4{loc_sram_buff_w15[158][4]}} & loc_sram_buff_w15[158][3:0]);
	loc_rdata_buff[ 387: 384] = ({4{loc_sram_buff_w0[159][4]}} & loc_sram_buff_w0[159][3:0]) | ({4{loc_sram_buff_w1[159][4]}} & loc_sram_buff_w1[159][3:0]) | ({4{loc_sram_buff_w2[159][4]}} & loc_sram_buff_w2[159][3:0]) | ({4{loc_sram_buff_w3[159][4]}} & loc_sram_buff_w3[159][3:0]) | ({4{loc_sram_buff_w4[159][4]}} & loc_sram_buff_w4[159][3:0]) | ({4{loc_sram_buff_w5[159][4]}} & loc_sram_buff_w5[159][3:0]) | ({4{loc_sram_buff_w6[159][4]}} & loc_sram_buff_w6[159][3:0]) | ({4{loc_sram_buff_w7[159][4]}} & loc_sram_buff_w7[159][3:0]) | ({4{loc_sram_buff_w8[159][4]}} & loc_sram_buff_w8[159][3:0]) | ({4{loc_sram_buff_w9[159][4]}} & loc_sram_buff_w9[159][3:0]) | ({4{loc_sram_buff_w10[159][4]}} & loc_sram_buff_w10[159][3:0]) | ({4{loc_sram_buff_w11[159][4]}} & loc_sram_buff_w11[159][3:0]) | ({4{loc_sram_buff_w12[159][4]}} & loc_sram_buff_w12[159][3:0]) | ({4{loc_sram_buff_w13[159][4]}} & loc_sram_buff_w13[159][3:0]) | ({4{loc_sram_buff_w14[159][4]}} & loc_sram_buff_w14[159][3:0]) | ({4{loc_sram_buff_w15[159][4]}} & loc_sram_buff_w15[159][3:0]);
	loc_rdata_buff[ 383: 380] = ({4{loc_sram_buff_w0[160][4]}} & loc_sram_buff_w0[160][3:0]) | ({4{loc_sram_buff_w1[160][4]}} & loc_sram_buff_w1[160][3:0]) | ({4{loc_sram_buff_w2[160][4]}} & loc_sram_buff_w2[160][3:0]) | ({4{loc_sram_buff_w3[160][4]}} & loc_sram_buff_w3[160][3:0]) | ({4{loc_sram_buff_w4[160][4]}} & loc_sram_buff_w4[160][3:0]) | ({4{loc_sram_buff_w5[160][4]}} & loc_sram_buff_w5[160][3:0]) | ({4{loc_sram_buff_w6[160][4]}} & loc_sram_buff_w6[160][3:0]) | ({4{loc_sram_buff_w7[160][4]}} & loc_sram_buff_w7[160][3:0]) | ({4{loc_sram_buff_w8[160][4]}} & loc_sram_buff_w8[160][3:0]) | ({4{loc_sram_buff_w9[160][4]}} & loc_sram_buff_w9[160][3:0]) | ({4{loc_sram_buff_w10[160][4]}} & loc_sram_buff_w10[160][3:0]) | ({4{loc_sram_buff_w11[160][4]}} & loc_sram_buff_w11[160][3:0]) | ({4{loc_sram_buff_w12[160][4]}} & loc_sram_buff_w12[160][3:0]) | ({4{loc_sram_buff_w13[160][4]}} & loc_sram_buff_w13[160][3:0]) | ({4{loc_sram_buff_w14[160][4]}} & loc_sram_buff_w14[160][3:0]) | ({4{loc_sram_buff_w15[160][4]}} & loc_sram_buff_w15[160][3:0]);
	loc_rdata_buff[ 379: 376] = ({4{loc_sram_buff_w0[161][4]}} & loc_sram_buff_w0[161][3:0]) | ({4{loc_sram_buff_w1[161][4]}} & loc_sram_buff_w1[161][3:0]) | ({4{loc_sram_buff_w2[161][4]}} & loc_sram_buff_w2[161][3:0]) | ({4{loc_sram_buff_w3[161][4]}} & loc_sram_buff_w3[161][3:0]) | ({4{loc_sram_buff_w4[161][4]}} & loc_sram_buff_w4[161][3:0]) | ({4{loc_sram_buff_w5[161][4]}} & loc_sram_buff_w5[161][3:0]) | ({4{loc_sram_buff_w6[161][4]}} & loc_sram_buff_w6[161][3:0]) | ({4{loc_sram_buff_w7[161][4]}} & loc_sram_buff_w7[161][3:0]) | ({4{loc_sram_buff_w8[161][4]}} & loc_sram_buff_w8[161][3:0]) | ({4{loc_sram_buff_w9[161][4]}} & loc_sram_buff_w9[161][3:0]) | ({4{loc_sram_buff_w10[161][4]}} & loc_sram_buff_w10[161][3:0]) | ({4{loc_sram_buff_w11[161][4]}} & loc_sram_buff_w11[161][3:0]) | ({4{loc_sram_buff_w12[161][4]}} & loc_sram_buff_w12[161][3:0]) | ({4{loc_sram_buff_w13[161][4]}} & loc_sram_buff_w13[161][3:0]) | ({4{loc_sram_buff_w14[161][4]}} & loc_sram_buff_w14[161][3:0]) | ({4{loc_sram_buff_w15[161][4]}} & loc_sram_buff_w15[161][3:0]);
	loc_rdata_buff[ 375: 372] = ({4{loc_sram_buff_w0[162][4]}} & loc_sram_buff_w0[162][3:0]) | ({4{loc_sram_buff_w1[162][4]}} & loc_sram_buff_w1[162][3:0]) | ({4{loc_sram_buff_w2[162][4]}} & loc_sram_buff_w2[162][3:0]) | ({4{loc_sram_buff_w3[162][4]}} & loc_sram_buff_w3[162][3:0]) | ({4{loc_sram_buff_w4[162][4]}} & loc_sram_buff_w4[162][3:0]) | ({4{loc_sram_buff_w5[162][4]}} & loc_sram_buff_w5[162][3:0]) | ({4{loc_sram_buff_w6[162][4]}} & loc_sram_buff_w6[162][3:0]) | ({4{loc_sram_buff_w7[162][4]}} & loc_sram_buff_w7[162][3:0]) | ({4{loc_sram_buff_w8[162][4]}} & loc_sram_buff_w8[162][3:0]) | ({4{loc_sram_buff_w9[162][4]}} & loc_sram_buff_w9[162][3:0]) | ({4{loc_sram_buff_w10[162][4]}} & loc_sram_buff_w10[162][3:0]) | ({4{loc_sram_buff_w11[162][4]}} & loc_sram_buff_w11[162][3:0]) | ({4{loc_sram_buff_w12[162][4]}} & loc_sram_buff_w12[162][3:0]) | ({4{loc_sram_buff_w13[162][4]}} & loc_sram_buff_w13[162][3:0]) | ({4{loc_sram_buff_w14[162][4]}} & loc_sram_buff_w14[162][3:0]) | ({4{loc_sram_buff_w15[162][4]}} & loc_sram_buff_w15[162][3:0]);
	loc_rdata_buff[ 371: 368] = ({4{loc_sram_buff_w0[163][4]}} & loc_sram_buff_w0[163][3:0]) | ({4{loc_sram_buff_w1[163][4]}} & loc_sram_buff_w1[163][3:0]) | ({4{loc_sram_buff_w2[163][4]}} & loc_sram_buff_w2[163][3:0]) | ({4{loc_sram_buff_w3[163][4]}} & loc_sram_buff_w3[163][3:0]) | ({4{loc_sram_buff_w4[163][4]}} & loc_sram_buff_w4[163][3:0]) | ({4{loc_sram_buff_w5[163][4]}} & loc_sram_buff_w5[163][3:0]) | ({4{loc_sram_buff_w6[163][4]}} & loc_sram_buff_w6[163][3:0]) | ({4{loc_sram_buff_w7[163][4]}} & loc_sram_buff_w7[163][3:0]) | ({4{loc_sram_buff_w8[163][4]}} & loc_sram_buff_w8[163][3:0]) | ({4{loc_sram_buff_w9[163][4]}} & loc_sram_buff_w9[163][3:0]) | ({4{loc_sram_buff_w10[163][4]}} & loc_sram_buff_w10[163][3:0]) | ({4{loc_sram_buff_w11[163][4]}} & loc_sram_buff_w11[163][3:0]) | ({4{loc_sram_buff_w12[163][4]}} & loc_sram_buff_w12[163][3:0]) | ({4{loc_sram_buff_w13[163][4]}} & loc_sram_buff_w13[163][3:0]) | ({4{loc_sram_buff_w14[163][4]}} & loc_sram_buff_w14[163][3:0]) | ({4{loc_sram_buff_w15[163][4]}} & loc_sram_buff_w15[163][3:0]);
	loc_rdata_buff[ 367: 364] = ({4{loc_sram_buff_w0[164][4]}} & loc_sram_buff_w0[164][3:0]) | ({4{loc_sram_buff_w1[164][4]}} & loc_sram_buff_w1[164][3:0]) | ({4{loc_sram_buff_w2[164][4]}} & loc_sram_buff_w2[164][3:0]) | ({4{loc_sram_buff_w3[164][4]}} & loc_sram_buff_w3[164][3:0]) | ({4{loc_sram_buff_w4[164][4]}} & loc_sram_buff_w4[164][3:0]) | ({4{loc_sram_buff_w5[164][4]}} & loc_sram_buff_w5[164][3:0]) | ({4{loc_sram_buff_w6[164][4]}} & loc_sram_buff_w6[164][3:0]) | ({4{loc_sram_buff_w7[164][4]}} & loc_sram_buff_w7[164][3:0]) | ({4{loc_sram_buff_w8[164][4]}} & loc_sram_buff_w8[164][3:0]) | ({4{loc_sram_buff_w9[164][4]}} & loc_sram_buff_w9[164][3:0]) | ({4{loc_sram_buff_w10[164][4]}} & loc_sram_buff_w10[164][3:0]) | ({4{loc_sram_buff_w11[164][4]}} & loc_sram_buff_w11[164][3:0]) | ({4{loc_sram_buff_w12[164][4]}} & loc_sram_buff_w12[164][3:0]) | ({4{loc_sram_buff_w13[164][4]}} & loc_sram_buff_w13[164][3:0]) | ({4{loc_sram_buff_w14[164][4]}} & loc_sram_buff_w14[164][3:0]) | ({4{loc_sram_buff_w15[164][4]}} & loc_sram_buff_w15[164][3:0]);
	loc_rdata_buff[ 363: 360] = ({4{loc_sram_buff_w0[165][4]}} & loc_sram_buff_w0[165][3:0]) | ({4{loc_sram_buff_w1[165][4]}} & loc_sram_buff_w1[165][3:0]) | ({4{loc_sram_buff_w2[165][4]}} & loc_sram_buff_w2[165][3:0]) | ({4{loc_sram_buff_w3[165][4]}} & loc_sram_buff_w3[165][3:0]) | ({4{loc_sram_buff_w4[165][4]}} & loc_sram_buff_w4[165][3:0]) | ({4{loc_sram_buff_w5[165][4]}} & loc_sram_buff_w5[165][3:0]) | ({4{loc_sram_buff_w6[165][4]}} & loc_sram_buff_w6[165][3:0]) | ({4{loc_sram_buff_w7[165][4]}} & loc_sram_buff_w7[165][3:0]) | ({4{loc_sram_buff_w8[165][4]}} & loc_sram_buff_w8[165][3:0]) | ({4{loc_sram_buff_w9[165][4]}} & loc_sram_buff_w9[165][3:0]) | ({4{loc_sram_buff_w10[165][4]}} & loc_sram_buff_w10[165][3:0]) | ({4{loc_sram_buff_w11[165][4]}} & loc_sram_buff_w11[165][3:0]) | ({4{loc_sram_buff_w12[165][4]}} & loc_sram_buff_w12[165][3:0]) | ({4{loc_sram_buff_w13[165][4]}} & loc_sram_buff_w13[165][3:0]) | ({4{loc_sram_buff_w14[165][4]}} & loc_sram_buff_w14[165][3:0]) | ({4{loc_sram_buff_w15[165][4]}} & loc_sram_buff_w15[165][3:0]);
	loc_rdata_buff[ 359: 356] = ({4{loc_sram_buff_w0[166][4]}} & loc_sram_buff_w0[166][3:0]) | ({4{loc_sram_buff_w1[166][4]}} & loc_sram_buff_w1[166][3:0]) | ({4{loc_sram_buff_w2[166][4]}} & loc_sram_buff_w2[166][3:0]) | ({4{loc_sram_buff_w3[166][4]}} & loc_sram_buff_w3[166][3:0]) | ({4{loc_sram_buff_w4[166][4]}} & loc_sram_buff_w4[166][3:0]) | ({4{loc_sram_buff_w5[166][4]}} & loc_sram_buff_w5[166][3:0]) | ({4{loc_sram_buff_w6[166][4]}} & loc_sram_buff_w6[166][3:0]) | ({4{loc_sram_buff_w7[166][4]}} & loc_sram_buff_w7[166][3:0]) | ({4{loc_sram_buff_w8[166][4]}} & loc_sram_buff_w8[166][3:0]) | ({4{loc_sram_buff_w9[166][4]}} & loc_sram_buff_w9[166][3:0]) | ({4{loc_sram_buff_w10[166][4]}} & loc_sram_buff_w10[166][3:0]) | ({4{loc_sram_buff_w11[166][4]}} & loc_sram_buff_w11[166][3:0]) | ({4{loc_sram_buff_w12[166][4]}} & loc_sram_buff_w12[166][3:0]) | ({4{loc_sram_buff_w13[166][4]}} & loc_sram_buff_w13[166][3:0]) | ({4{loc_sram_buff_w14[166][4]}} & loc_sram_buff_w14[166][3:0]) | ({4{loc_sram_buff_w15[166][4]}} & loc_sram_buff_w15[166][3:0]);
	loc_rdata_buff[ 355: 352] = ({4{loc_sram_buff_w0[167][4]}} & loc_sram_buff_w0[167][3:0]) | ({4{loc_sram_buff_w1[167][4]}} & loc_sram_buff_w1[167][3:0]) | ({4{loc_sram_buff_w2[167][4]}} & loc_sram_buff_w2[167][3:0]) | ({4{loc_sram_buff_w3[167][4]}} & loc_sram_buff_w3[167][3:0]) | ({4{loc_sram_buff_w4[167][4]}} & loc_sram_buff_w4[167][3:0]) | ({4{loc_sram_buff_w5[167][4]}} & loc_sram_buff_w5[167][3:0]) | ({4{loc_sram_buff_w6[167][4]}} & loc_sram_buff_w6[167][3:0]) | ({4{loc_sram_buff_w7[167][4]}} & loc_sram_buff_w7[167][3:0]) | ({4{loc_sram_buff_w8[167][4]}} & loc_sram_buff_w8[167][3:0]) | ({4{loc_sram_buff_w9[167][4]}} & loc_sram_buff_w9[167][3:0]) | ({4{loc_sram_buff_w10[167][4]}} & loc_sram_buff_w10[167][3:0]) | ({4{loc_sram_buff_w11[167][4]}} & loc_sram_buff_w11[167][3:0]) | ({4{loc_sram_buff_w12[167][4]}} & loc_sram_buff_w12[167][3:0]) | ({4{loc_sram_buff_w13[167][4]}} & loc_sram_buff_w13[167][3:0]) | ({4{loc_sram_buff_w14[167][4]}} & loc_sram_buff_w14[167][3:0]) | ({4{loc_sram_buff_w15[167][4]}} & loc_sram_buff_w15[167][3:0]);
	loc_rdata_buff[ 351: 348] = ({4{loc_sram_buff_w0[168][4]}} & loc_sram_buff_w0[168][3:0]) | ({4{loc_sram_buff_w1[168][4]}} & loc_sram_buff_w1[168][3:0]) | ({4{loc_sram_buff_w2[168][4]}} & loc_sram_buff_w2[168][3:0]) | ({4{loc_sram_buff_w3[168][4]}} & loc_sram_buff_w3[168][3:0]) | ({4{loc_sram_buff_w4[168][4]}} & loc_sram_buff_w4[168][3:0]) | ({4{loc_sram_buff_w5[168][4]}} & loc_sram_buff_w5[168][3:0]) | ({4{loc_sram_buff_w6[168][4]}} & loc_sram_buff_w6[168][3:0]) | ({4{loc_sram_buff_w7[168][4]}} & loc_sram_buff_w7[168][3:0]) | ({4{loc_sram_buff_w8[168][4]}} & loc_sram_buff_w8[168][3:0]) | ({4{loc_sram_buff_w9[168][4]}} & loc_sram_buff_w9[168][3:0]) | ({4{loc_sram_buff_w10[168][4]}} & loc_sram_buff_w10[168][3:0]) | ({4{loc_sram_buff_w11[168][4]}} & loc_sram_buff_w11[168][3:0]) | ({4{loc_sram_buff_w12[168][4]}} & loc_sram_buff_w12[168][3:0]) | ({4{loc_sram_buff_w13[168][4]}} & loc_sram_buff_w13[168][3:0]) | ({4{loc_sram_buff_w14[168][4]}} & loc_sram_buff_w14[168][3:0]) | ({4{loc_sram_buff_w15[168][4]}} & loc_sram_buff_w15[168][3:0]);
	loc_rdata_buff[ 347: 344] = ({4{loc_sram_buff_w0[169][4]}} & loc_sram_buff_w0[169][3:0]) | ({4{loc_sram_buff_w1[169][4]}} & loc_sram_buff_w1[169][3:0]) | ({4{loc_sram_buff_w2[169][4]}} & loc_sram_buff_w2[169][3:0]) | ({4{loc_sram_buff_w3[169][4]}} & loc_sram_buff_w3[169][3:0]) | ({4{loc_sram_buff_w4[169][4]}} & loc_sram_buff_w4[169][3:0]) | ({4{loc_sram_buff_w5[169][4]}} & loc_sram_buff_w5[169][3:0]) | ({4{loc_sram_buff_w6[169][4]}} & loc_sram_buff_w6[169][3:0]) | ({4{loc_sram_buff_w7[169][4]}} & loc_sram_buff_w7[169][3:0]) | ({4{loc_sram_buff_w8[169][4]}} & loc_sram_buff_w8[169][3:0]) | ({4{loc_sram_buff_w9[169][4]}} & loc_sram_buff_w9[169][3:0]) | ({4{loc_sram_buff_w10[169][4]}} & loc_sram_buff_w10[169][3:0]) | ({4{loc_sram_buff_w11[169][4]}} & loc_sram_buff_w11[169][3:0]) | ({4{loc_sram_buff_w12[169][4]}} & loc_sram_buff_w12[169][3:0]) | ({4{loc_sram_buff_w13[169][4]}} & loc_sram_buff_w13[169][3:0]) | ({4{loc_sram_buff_w14[169][4]}} & loc_sram_buff_w14[169][3:0]) | ({4{loc_sram_buff_w15[169][4]}} & loc_sram_buff_w15[169][3:0]);
	loc_rdata_buff[ 343: 340] = ({4{loc_sram_buff_w0[170][4]}} & loc_sram_buff_w0[170][3:0]) | ({4{loc_sram_buff_w1[170][4]}} & loc_sram_buff_w1[170][3:0]) | ({4{loc_sram_buff_w2[170][4]}} & loc_sram_buff_w2[170][3:0]) | ({4{loc_sram_buff_w3[170][4]}} & loc_sram_buff_w3[170][3:0]) | ({4{loc_sram_buff_w4[170][4]}} & loc_sram_buff_w4[170][3:0]) | ({4{loc_sram_buff_w5[170][4]}} & loc_sram_buff_w5[170][3:0]) | ({4{loc_sram_buff_w6[170][4]}} & loc_sram_buff_w6[170][3:0]) | ({4{loc_sram_buff_w7[170][4]}} & loc_sram_buff_w7[170][3:0]) | ({4{loc_sram_buff_w8[170][4]}} & loc_sram_buff_w8[170][3:0]) | ({4{loc_sram_buff_w9[170][4]}} & loc_sram_buff_w9[170][3:0]) | ({4{loc_sram_buff_w10[170][4]}} & loc_sram_buff_w10[170][3:0]) | ({4{loc_sram_buff_w11[170][4]}} & loc_sram_buff_w11[170][3:0]) | ({4{loc_sram_buff_w12[170][4]}} & loc_sram_buff_w12[170][3:0]) | ({4{loc_sram_buff_w13[170][4]}} & loc_sram_buff_w13[170][3:0]) | ({4{loc_sram_buff_w14[170][4]}} & loc_sram_buff_w14[170][3:0]) | ({4{loc_sram_buff_w15[170][4]}} & loc_sram_buff_w15[170][3:0]);
	loc_rdata_buff[ 339: 336] = ({4{loc_sram_buff_w0[171][4]}} & loc_sram_buff_w0[171][3:0]) | ({4{loc_sram_buff_w1[171][4]}} & loc_sram_buff_w1[171][3:0]) | ({4{loc_sram_buff_w2[171][4]}} & loc_sram_buff_w2[171][3:0]) | ({4{loc_sram_buff_w3[171][4]}} & loc_sram_buff_w3[171][3:0]) | ({4{loc_sram_buff_w4[171][4]}} & loc_sram_buff_w4[171][3:0]) | ({4{loc_sram_buff_w5[171][4]}} & loc_sram_buff_w5[171][3:0]) | ({4{loc_sram_buff_w6[171][4]}} & loc_sram_buff_w6[171][3:0]) | ({4{loc_sram_buff_w7[171][4]}} & loc_sram_buff_w7[171][3:0]) | ({4{loc_sram_buff_w8[171][4]}} & loc_sram_buff_w8[171][3:0]) | ({4{loc_sram_buff_w9[171][4]}} & loc_sram_buff_w9[171][3:0]) | ({4{loc_sram_buff_w10[171][4]}} & loc_sram_buff_w10[171][3:0]) | ({4{loc_sram_buff_w11[171][4]}} & loc_sram_buff_w11[171][3:0]) | ({4{loc_sram_buff_w12[171][4]}} & loc_sram_buff_w12[171][3:0]) | ({4{loc_sram_buff_w13[171][4]}} & loc_sram_buff_w13[171][3:0]) | ({4{loc_sram_buff_w14[171][4]}} & loc_sram_buff_w14[171][3:0]) | ({4{loc_sram_buff_w15[171][4]}} & loc_sram_buff_w15[171][3:0]);
	loc_rdata_buff[ 335: 332] = ({4{loc_sram_buff_w0[172][4]}} & loc_sram_buff_w0[172][3:0]) | ({4{loc_sram_buff_w1[172][4]}} & loc_sram_buff_w1[172][3:0]) | ({4{loc_sram_buff_w2[172][4]}} & loc_sram_buff_w2[172][3:0]) | ({4{loc_sram_buff_w3[172][4]}} & loc_sram_buff_w3[172][3:0]) | ({4{loc_sram_buff_w4[172][4]}} & loc_sram_buff_w4[172][3:0]) | ({4{loc_sram_buff_w5[172][4]}} & loc_sram_buff_w5[172][3:0]) | ({4{loc_sram_buff_w6[172][4]}} & loc_sram_buff_w6[172][3:0]) | ({4{loc_sram_buff_w7[172][4]}} & loc_sram_buff_w7[172][3:0]) | ({4{loc_sram_buff_w8[172][4]}} & loc_sram_buff_w8[172][3:0]) | ({4{loc_sram_buff_w9[172][4]}} & loc_sram_buff_w9[172][3:0]) | ({4{loc_sram_buff_w10[172][4]}} & loc_sram_buff_w10[172][3:0]) | ({4{loc_sram_buff_w11[172][4]}} & loc_sram_buff_w11[172][3:0]) | ({4{loc_sram_buff_w12[172][4]}} & loc_sram_buff_w12[172][3:0]) | ({4{loc_sram_buff_w13[172][4]}} & loc_sram_buff_w13[172][3:0]) | ({4{loc_sram_buff_w14[172][4]}} & loc_sram_buff_w14[172][3:0]) | ({4{loc_sram_buff_w15[172][4]}} & loc_sram_buff_w15[172][3:0]);
	loc_rdata_buff[ 331: 328] = ({4{loc_sram_buff_w0[173][4]}} & loc_sram_buff_w0[173][3:0]) | ({4{loc_sram_buff_w1[173][4]}} & loc_sram_buff_w1[173][3:0]) | ({4{loc_sram_buff_w2[173][4]}} & loc_sram_buff_w2[173][3:0]) | ({4{loc_sram_buff_w3[173][4]}} & loc_sram_buff_w3[173][3:0]) | ({4{loc_sram_buff_w4[173][4]}} & loc_sram_buff_w4[173][3:0]) | ({4{loc_sram_buff_w5[173][4]}} & loc_sram_buff_w5[173][3:0]) | ({4{loc_sram_buff_w6[173][4]}} & loc_sram_buff_w6[173][3:0]) | ({4{loc_sram_buff_w7[173][4]}} & loc_sram_buff_w7[173][3:0]) | ({4{loc_sram_buff_w8[173][4]}} & loc_sram_buff_w8[173][3:0]) | ({4{loc_sram_buff_w9[173][4]}} & loc_sram_buff_w9[173][3:0]) | ({4{loc_sram_buff_w10[173][4]}} & loc_sram_buff_w10[173][3:0]) | ({4{loc_sram_buff_w11[173][4]}} & loc_sram_buff_w11[173][3:0]) | ({4{loc_sram_buff_w12[173][4]}} & loc_sram_buff_w12[173][3:0]) | ({4{loc_sram_buff_w13[173][4]}} & loc_sram_buff_w13[173][3:0]) | ({4{loc_sram_buff_w14[173][4]}} & loc_sram_buff_w14[173][3:0]) | ({4{loc_sram_buff_w15[173][4]}} & loc_sram_buff_w15[173][3:0]);
	loc_rdata_buff[ 327: 324] = ({4{loc_sram_buff_w0[174][4]}} & loc_sram_buff_w0[174][3:0]) | ({4{loc_sram_buff_w1[174][4]}} & loc_sram_buff_w1[174][3:0]) | ({4{loc_sram_buff_w2[174][4]}} & loc_sram_buff_w2[174][3:0]) | ({4{loc_sram_buff_w3[174][4]}} & loc_sram_buff_w3[174][3:0]) | ({4{loc_sram_buff_w4[174][4]}} & loc_sram_buff_w4[174][3:0]) | ({4{loc_sram_buff_w5[174][4]}} & loc_sram_buff_w5[174][3:0]) | ({4{loc_sram_buff_w6[174][4]}} & loc_sram_buff_w6[174][3:0]) | ({4{loc_sram_buff_w7[174][4]}} & loc_sram_buff_w7[174][3:0]) | ({4{loc_sram_buff_w8[174][4]}} & loc_sram_buff_w8[174][3:0]) | ({4{loc_sram_buff_w9[174][4]}} & loc_sram_buff_w9[174][3:0]) | ({4{loc_sram_buff_w10[174][4]}} & loc_sram_buff_w10[174][3:0]) | ({4{loc_sram_buff_w11[174][4]}} & loc_sram_buff_w11[174][3:0]) | ({4{loc_sram_buff_w12[174][4]}} & loc_sram_buff_w12[174][3:0]) | ({4{loc_sram_buff_w13[174][4]}} & loc_sram_buff_w13[174][3:0]) | ({4{loc_sram_buff_w14[174][4]}} & loc_sram_buff_w14[174][3:0]) | ({4{loc_sram_buff_w15[174][4]}} & loc_sram_buff_w15[174][3:0]);
	loc_rdata_buff[ 323: 320] = ({4{loc_sram_buff_w0[175][4]}} & loc_sram_buff_w0[175][3:0]) | ({4{loc_sram_buff_w1[175][4]}} & loc_sram_buff_w1[175][3:0]) | ({4{loc_sram_buff_w2[175][4]}} & loc_sram_buff_w2[175][3:0]) | ({4{loc_sram_buff_w3[175][4]}} & loc_sram_buff_w3[175][3:0]) | ({4{loc_sram_buff_w4[175][4]}} & loc_sram_buff_w4[175][3:0]) | ({4{loc_sram_buff_w5[175][4]}} & loc_sram_buff_w5[175][3:0]) | ({4{loc_sram_buff_w6[175][4]}} & loc_sram_buff_w6[175][3:0]) | ({4{loc_sram_buff_w7[175][4]}} & loc_sram_buff_w7[175][3:0]) | ({4{loc_sram_buff_w8[175][4]}} & loc_sram_buff_w8[175][3:0]) | ({4{loc_sram_buff_w9[175][4]}} & loc_sram_buff_w9[175][3:0]) | ({4{loc_sram_buff_w10[175][4]}} & loc_sram_buff_w10[175][3:0]) | ({4{loc_sram_buff_w11[175][4]}} & loc_sram_buff_w11[175][3:0]) | ({4{loc_sram_buff_w12[175][4]}} & loc_sram_buff_w12[175][3:0]) | ({4{loc_sram_buff_w13[175][4]}} & loc_sram_buff_w13[175][3:0]) | ({4{loc_sram_buff_w14[175][4]}} & loc_sram_buff_w14[175][3:0]) | ({4{loc_sram_buff_w15[175][4]}} & loc_sram_buff_w15[175][3:0]);
	loc_rdata_buff[ 319: 316] = ({4{loc_sram_buff_w0[176][4]}} & loc_sram_buff_w0[176][3:0]) | ({4{loc_sram_buff_w1[176][4]}} & loc_sram_buff_w1[176][3:0]) | ({4{loc_sram_buff_w2[176][4]}} & loc_sram_buff_w2[176][3:0]) | ({4{loc_sram_buff_w3[176][4]}} & loc_sram_buff_w3[176][3:0]) | ({4{loc_sram_buff_w4[176][4]}} & loc_sram_buff_w4[176][3:0]) | ({4{loc_sram_buff_w5[176][4]}} & loc_sram_buff_w5[176][3:0]) | ({4{loc_sram_buff_w6[176][4]}} & loc_sram_buff_w6[176][3:0]) | ({4{loc_sram_buff_w7[176][4]}} & loc_sram_buff_w7[176][3:0]) | ({4{loc_sram_buff_w8[176][4]}} & loc_sram_buff_w8[176][3:0]) | ({4{loc_sram_buff_w9[176][4]}} & loc_sram_buff_w9[176][3:0]) | ({4{loc_sram_buff_w10[176][4]}} & loc_sram_buff_w10[176][3:0]) | ({4{loc_sram_buff_w11[176][4]}} & loc_sram_buff_w11[176][3:0]) | ({4{loc_sram_buff_w12[176][4]}} & loc_sram_buff_w12[176][3:0]) | ({4{loc_sram_buff_w13[176][4]}} & loc_sram_buff_w13[176][3:0]) | ({4{loc_sram_buff_w14[176][4]}} & loc_sram_buff_w14[176][3:0]) | ({4{loc_sram_buff_w15[176][4]}} & loc_sram_buff_w15[176][3:0]);
	loc_rdata_buff[ 315: 312] = ({4{loc_sram_buff_w0[177][4]}} & loc_sram_buff_w0[177][3:0]) | ({4{loc_sram_buff_w1[177][4]}} & loc_sram_buff_w1[177][3:0]) | ({4{loc_sram_buff_w2[177][4]}} & loc_sram_buff_w2[177][3:0]) | ({4{loc_sram_buff_w3[177][4]}} & loc_sram_buff_w3[177][3:0]) | ({4{loc_sram_buff_w4[177][4]}} & loc_sram_buff_w4[177][3:0]) | ({4{loc_sram_buff_w5[177][4]}} & loc_sram_buff_w5[177][3:0]) | ({4{loc_sram_buff_w6[177][4]}} & loc_sram_buff_w6[177][3:0]) | ({4{loc_sram_buff_w7[177][4]}} & loc_sram_buff_w7[177][3:0]) | ({4{loc_sram_buff_w8[177][4]}} & loc_sram_buff_w8[177][3:0]) | ({4{loc_sram_buff_w9[177][4]}} & loc_sram_buff_w9[177][3:0]) | ({4{loc_sram_buff_w10[177][4]}} & loc_sram_buff_w10[177][3:0]) | ({4{loc_sram_buff_w11[177][4]}} & loc_sram_buff_w11[177][3:0]) | ({4{loc_sram_buff_w12[177][4]}} & loc_sram_buff_w12[177][3:0]) | ({4{loc_sram_buff_w13[177][4]}} & loc_sram_buff_w13[177][3:0]) | ({4{loc_sram_buff_w14[177][4]}} & loc_sram_buff_w14[177][3:0]) | ({4{loc_sram_buff_w15[177][4]}} & loc_sram_buff_w15[177][3:0]);
	loc_rdata_buff[ 311: 308] = ({4{loc_sram_buff_w0[178][4]}} & loc_sram_buff_w0[178][3:0]) | ({4{loc_sram_buff_w1[178][4]}} & loc_sram_buff_w1[178][3:0]) | ({4{loc_sram_buff_w2[178][4]}} & loc_sram_buff_w2[178][3:0]) | ({4{loc_sram_buff_w3[178][4]}} & loc_sram_buff_w3[178][3:0]) | ({4{loc_sram_buff_w4[178][4]}} & loc_sram_buff_w4[178][3:0]) | ({4{loc_sram_buff_w5[178][4]}} & loc_sram_buff_w5[178][3:0]) | ({4{loc_sram_buff_w6[178][4]}} & loc_sram_buff_w6[178][3:0]) | ({4{loc_sram_buff_w7[178][4]}} & loc_sram_buff_w7[178][3:0]) | ({4{loc_sram_buff_w8[178][4]}} & loc_sram_buff_w8[178][3:0]) | ({4{loc_sram_buff_w9[178][4]}} & loc_sram_buff_w9[178][3:0]) | ({4{loc_sram_buff_w10[178][4]}} & loc_sram_buff_w10[178][3:0]) | ({4{loc_sram_buff_w11[178][4]}} & loc_sram_buff_w11[178][3:0]) | ({4{loc_sram_buff_w12[178][4]}} & loc_sram_buff_w12[178][3:0]) | ({4{loc_sram_buff_w13[178][4]}} & loc_sram_buff_w13[178][3:0]) | ({4{loc_sram_buff_w14[178][4]}} & loc_sram_buff_w14[178][3:0]) | ({4{loc_sram_buff_w15[178][4]}} & loc_sram_buff_w15[178][3:0]);
	loc_rdata_buff[ 307: 304] = ({4{loc_sram_buff_w0[179][4]}} & loc_sram_buff_w0[179][3:0]) | ({4{loc_sram_buff_w1[179][4]}} & loc_sram_buff_w1[179][3:0]) | ({4{loc_sram_buff_w2[179][4]}} & loc_sram_buff_w2[179][3:0]) | ({4{loc_sram_buff_w3[179][4]}} & loc_sram_buff_w3[179][3:0]) | ({4{loc_sram_buff_w4[179][4]}} & loc_sram_buff_w4[179][3:0]) | ({4{loc_sram_buff_w5[179][4]}} & loc_sram_buff_w5[179][3:0]) | ({4{loc_sram_buff_w6[179][4]}} & loc_sram_buff_w6[179][3:0]) | ({4{loc_sram_buff_w7[179][4]}} & loc_sram_buff_w7[179][3:0]) | ({4{loc_sram_buff_w8[179][4]}} & loc_sram_buff_w8[179][3:0]) | ({4{loc_sram_buff_w9[179][4]}} & loc_sram_buff_w9[179][3:0]) | ({4{loc_sram_buff_w10[179][4]}} & loc_sram_buff_w10[179][3:0]) | ({4{loc_sram_buff_w11[179][4]}} & loc_sram_buff_w11[179][3:0]) | ({4{loc_sram_buff_w12[179][4]}} & loc_sram_buff_w12[179][3:0]) | ({4{loc_sram_buff_w13[179][4]}} & loc_sram_buff_w13[179][3:0]) | ({4{loc_sram_buff_w14[179][4]}} & loc_sram_buff_w14[179][3:0]) | ({4{loc_sram_buff_w15[179][4]}} & loc_sram_buff_w15[179][3:0]);
	loc_rdata_buff[ 303: 300] = ({4{loc_sram_buff_w0[180][4]}} & loc_sram_buff_w0[180][3:0]) | ({4{loc_sram_buff_w1[180][4]}} & loc_sram_buff_w1[180][3:0]) | ({4{loc_sram_buff_w2[180][4]}} & loc_sram_buff_w2[180][3:0]) | ({4{loc_sram_buff_w3[180][4]}} & loc_sram_buff_w3[180][3:0]) | ({4{loc_sram_buff_w4[180][4]}} & loc_sram_buff_w4[180][3:0]) | ({4{loc_sram_buff_w5[180][4]}} & loc_sram_buff_w5[180][3:0]) | ({4{loc_sram_buff_w6[180][4]}} & loc_sram_buff_w6[180][3:0]) | ({4{loc_sram_buff_w7[180][4]}} & loc_sram_buff_w7[180][3:0]) | ({4{loc_sram_buff_w8[180][4]}} & loc_sram_buff_w8[180][3:0]) | ({4{loc_sram_buff_w9[180][4]}} & loc_sram_buff_w9[180][3:0]) | ({4{loc_sram_buff_w10[180][4]}} & loc_sram_buff_w10[180][3:0]) | ({4{loc_sram_buff_w11[180][4]}} & loc_sram_buff_w11[180][3:0]) | ({4{loc_sram_buff_w12[180][4]}} & loc_sram_buff_w12[180][3:0]) | ({4{loc_sram_buff_w13[180][4]}} & loc_sram_buff_w13[180][3:0]) | ({4{loc_sram_buff_w14[180][4]}} & loc_sram_buff_w14[180][3:0]) | ({4{loc_sram_buff_w15[180][4]}} & loc_sram_buff_w15[180][3:0]);
	loc_rdata_buff[ 299: 296] = ({4{loc_sram_buff_w0[181][4]}} & loc_sram_buff_w0[181][3:0]) | ({4{loc_sram_buff_w1[181][4]}} & loc_sram_buff_w1[181][3:0]) | ({4{loc_sram_buff_w2[181][4]}} & loc_sram_buff_w2[181][3:0]) | ({4{loc_sram_buff_w3[181][4]}} & loc_sram_buff_w3[181][3:0]) | ({4{loc_sram_buff_w4[181][4]}} & loc_sram_buff_w4[181][3:0]) | ({4{loc_sram_buff_w5[181][4]}} & loc_sram_buff_w5[181][3:0]) | ({4{loc_sram_buff_w6[181][4]}} & loc_sram_buff_w6[181][3:0]) | ({4{loc_sram_buff_w7[181][4]}} & loc_sram_buff_w7[181][3:0]) | ({4{loc_sram_buff_w8[181][4]}} & loc_sram_buff_w8[181][3:0]) | ({4{loc_sram_buff_w9[181][4]}} & loc_sram_buff_w9[181][3:0]) | ({4{loc_sram_buff_w10[181][4]}} & loc_sram_buff_w10[181][3:0]) | ({4{loc_sram_buff_w11[181][4]}} & loc_sram_buff_w11[181][3:0]) | ({4{loc_sram_buff_w12[181][4]}} & loc_sram_buff_w12[181][3:0]) | ({4{loc_sram_buff_w13[181][4]}} & loc_sram_buff_w13[181][3:0]) | ({4{loc_sram_buff_w14[181][4]}} & loc_sram_buff_w14[181][3:0]) | ({4{loc_sram_buff_w15[181][4]}} & loc_sram_buff_w15[181][3:0]);
	loc_rdata_buff[ 295: 292] = ({4{loc_sram_buff_w0[182][4]}} & loc_sram_buff_w0[182][3:0]) | ({4{loc_sram_buff_w1[182][4]}} & loc_sram_buff_w1[182][3:0]) | ({4{loc_sram_buff_w2[182][4]}} & loc_sram_buff_w2[182][3:0]) | ({4{loc_sram_buff_w3[182][4]}} & loc_sram_buff_w3[182][3:0]) | ({4{loc_sram_buff_w4[182][4]}} & loc_sram_buff_w4[182][3:0]) | ({4{loc_sram_buff_w5[182][4]}} & loc_sram_buff_w5[182][3:0]) | ({4{loc_sram_buff_w6[182][4]}} & loc_sram_buff_w6[182][3:0]) | ({4{loc_sram_buff_w7[182][4]}} & loc_sram_buff_w7[182][3:0]) | ({4{loc_sram_buff_w8[182][4]}} & loc_sram_buff_w8[182][3:0]) | ({4{loc_sram_buff_w9[182][4]}} & loc_sram_buff_w9[182][3:0]) | ({4{loc_sram_buff_w10[182][4]}} & loc_sram_buff_w10[182][3:0]) | ({4{loc_sram_buff_w11[182][4]}} & loc_sram_buff_w11[182][3:0]) | ({4{loc_sram_buff_w12[182][4]}} & loc_sram_buff_w12[182][3:0]) | ({4{loc_sram_buff_w13[182][4]}} & loc_sram_buff_w13[182][3:0]) | ({4{loc_sram_buff_w14[182][4]}} & loc_sram_buff_w14[182][3:0]) | ({4{loc_sram_buff_w15[182][4]}} & loc_sram_buff_w15[182][3:0]);
	loc_rdata_buff[ 291: 288] = ({4{loc_sram_buff_w0[183][4]}} & loc_sram_buff_w0[183][3:0]) | ({4{loc_sram_buff_w1[183][4]}} & loc_sram_buff_w1[183][3:0]) | ({4{loc_sram_buff_w2[183][4]}} & loc_sram_buff_w2[183][3:0]) | ({4{loc_sram_buff_w3[183][4]}} & loc_sram_buff_w3[183][3:0]) | ({4{loc_sram_buff_w4[183][4]}} & loc_sram_buff_w4[183][3:0]) | ({4{loc_sram_buff_w5[183][4]}} & loc_sram_buff_w5[183][3:0]) | ({4{loc_sram_buff_w6[183][4]}} & loc_sram_buff_w6[183][3:0]) | ({4{loc_sram_buff_w7[183][4]}} & loc_sram_buff_w7[183][3:0]) | ({4{loc_sram_buff_w8[183][4]}} & loc_sram_buff_w8[183][3:0]) | ({4{loc_sram_buff_w9[183][4]}} & loc_sram_buff_w9[183][3:0]) | ({4{loc_sram_buff_w10[183][4]}} & loc_sram_buff_w10[183][3:0]) | ({4{loc_sram_buff_w11[183][4]}} & loc_sram_buff_w11[183][3:0]) | ({4{loc_sram_buff_w12[183][4]}} & loc_sram_buff_w12[183][3:0]) | ({4{loc_sram_buff_w13[183][4]}} & loc_sram_buff_w13[183][3:0]) | ({4{loc_sram_buff_w14[183][4]}} & loc_sram_buff_w14[183][3:0]) | ({4{loc_sram_buff_w15[183][4]}} & loc_sram_buff_w15[183][3:0]);
	loc_rdata_buff[ 287: 284] = ({4{loc_sram_buff_w0[184][4]}} & loc_sram_buff_w0[184][3:0]) | ({4{loc_sram_buff_w1[184][4]}} & loc_sram_buff_w1[184][3:0]) | ({4{loc_sram_buff_w2[184][4]}} & loc_sram_buff_w2[184][3:0]) | ({4{loc_sram_buff_w3[184][4]}} & loc_sram_buff_w3[184][3:0]) | ({4{loc_sram_buff_w4[184][4]}} & loc_sram_buff_w4[184][3:0]) | ({4{loc_sram_buff_w5[184][4]}} & loc_sram_buff_w5[184][3:0]) | ({4{loc_sram_buff_w6[184][4]}} & loc_sram_buff_w6[184][3:0]) | ({4{loc_sram_buff_w7[184][4]}} & loc_sram_buff_w7[184][3:0]) | ({4{loc_sram_buff_w8[184][4]}} & loc_sram_buff_w8[184][3:0]) | ({4{loc_sram_buff_w9[184][4]}} & loc_sram_buff_w9[184][3:0]) | ({4{loc_sram_buff_w10[184][4]}} & loc_sram_buff_w10[184][3:0]) | ({4{loc_sram_buff_w11[184][4]}} & loc_sram_buff_w11[184][3:0]) | ({4{loc_sram_buff_w12[184][4]}} & loc_sram_buff_w12[184][3:0]) | ({4{loc_sram_buff_w13[184][4]}} & loc_sram_buff_w13[184][3:0]) | ({4{loc_sram_buff_w14[184][4]}} & loc_sram_buff_w14[184][3:0]) | ({4{loc_sram_buff_w15[184][4]}} & loc_sram_buff_w15[184][3:0]);
	loc_rdata_buff[ 283: 280] = ({4{loc_sram_buff_w0[185][4]}} & loc_sram_buff_w0[185][3:0]) | ({4{loc_sram_buff_w1[185][4]}} & loc_sram_buff_w1[185][3:0]) | ({4{loc_sram_buff_w2[185][4]}} & loc_sram_buff_w2[185][3:0]) | ({4{loc_sram_buff_w3[185][4]}} & loc_sram_buff_w3[185][3:0]) | ({4{loc_sram_buff_w4[185][4]}} & loc_sram_buff_w4[185][3:0]) | ({4{loc_sram_buff_w5[185][4]}} & loc_sram_buff_w5[185][3:0]) | ({4{loc_sram_buff_w6[185][4]}} & loc_sram_buff_w6[185][3:0]) | ({4{loc_sram_buff_w7[185][4]}} & loc_sram_buff_w7[185][3:0]) | ({4{loc_sram_buff_w8[185][4]}} & loc_sram_buff_w8[185][3:0]) | ({4{loc_sram_buff_w9[185][4]}} & loc_sram_buff_w9[185][3:0]) | ({4{loc_sram_buff_w10[185][4]}} & loc_sram_buff_w10[185][3:0]) | ({4{loc_sram_buff_w11[185][4]}} & loc_sram_buff_w11[185][3:0]) | ({4{loc_sram_buff_w12[185][4]}} & loc_sram_buff_w12[185][3:0]) | ({4{loc_sram_buff_w13[185][4]}} & loc_sram_buff_w13[185][3:0]) | ({4{loc_sram_buff_w14[185][4]}} & loc_sram_buff_w14[185][3:0]) | ({4{loc_sram_buff_w15[185][4]}} & loc_sram_buff_w15[185][3:0]);
	loc_rdata_buff[ 279: 276] = ({4{loc_sram_buff_w0[186][4]}} & loc_sram_buff_w0[186][3:0]) | ({4{loc_sram_buff_w1[186][4]}} & loc_sram_buff_w1[186][3:0]) | ({4{loc_sram_buff_w2[186][4]}} & loc_sram_buff_w2[186][3:0]) | ({4{loc_sram_buff_w3[186][4]}} & loc_sram_buff_w3[186][3:0]) | ({4{loc_sram_buff_w4[186][4]}} & loc_sram_buff_w4[186][3:0]) | ({4{loc_sram_buff_w5[186][4]}} & loc_sram_buff_w5[186][3:0]) | ({4{loc_sram_buff_w6[186][4]}} & loc_sram_buff_w6[186][3:0]) | ({4{loc_sram_buff_w7[186][4]}} & loc_sram_buff_w7[186][3:0]) | ({4{loc_sram_buff_w8[186][4]}} & loc_sram_buff_w8[186][3:0]) | ({4{loc_sram_buff_w9[186][4]}} & loc_sram_buff_w9[186][3:0]) | ({4{loc_sram_buff_w10[186][4]}} & loc_sram_buff_w10[186][3:0]) | ({4{loc_sram_buff_w11[186][4]}} & loc_sram_buff_w11[186][3:0]) | ({4{loc_sram_buff_w12[186][4]}} & loc_sram_buff_w12[186][3:0]) | ({4{loc_sram_buff_w13[186][4]}} & loc_sram_buff_w13[186][3:0]) | ({4{loc_sram_buff_w14[186][4]}} & loc_sram_buff_w14[186][3:0]) | ({4{loc_sram_buff_w15[186][4]}} & loc_sram_buff_w15[186][3:0]);
	loc_rdata_buff[ 275: 272] = ({4{loc_sram_buff_w0[187][4]}} & loc_sram_buff_w0[187][3:0]) | ({4{loc_sram_buff_w1[187][4]}} & loc_sram_buff_w1[187][3:0]) | ({4{loc_sram_buff_w2[187][4]}} & loc_sram_buff_w2[187][3:0]) | ({4{loc_sram_buff_w3[187][4]}} & loc_sram_buff_w3[187][3:0]) | ({4{loc_sram_buff_w4[187][4]}} & loc_sram_buff_w4[187][3:0]) | ({4{loc_sram_buff_w5[187][4]}} & loc_sram_buff_w5[187][3:0]) | ({4{loc_sram_buff_w6[187][4]}} & loc_sram_buff_w6[187][3:0]) | ({4{loc_sram_buff_w7[187][4]}} & loc_sram_buff_w7[187][3:0]) | ({4{loc_sram_buff_w8[187][4]}} & loc_sram_buff_w8[187][3:0]) | ({4{loc_sram_buff_w9[187][4]}} & loc_sram_buff_w9[187][3:0]) | ({4{loc_sram_buff_w10[187][4]}} & loc_sram_buff_w10[187][3:0]) | ({4{loc_sram_buff_w11[187][4]}} & loc_sram_buff_w11[187][3:0]) | ({4{loc_sram_buff_w12[187][4]}} & loc_sram_buff_w12[187][3:0]) | ({4{loc_sram_buff_w13[187][4]}} & loc_sram_buff_w13[187][3:0]) | ({4{loc_sram_buff_w14[187][4]}} & loc_sram_buff_w14[187][3:0]) | ({4{loc_sram_buff_w15[187][4]}} & loc_sram_buff_w15[187][3:0]);
	loc_rdata_buff[ 271: 268] = ({4{loc_sram_buff_w0[188][4]}} & loc_sram_buff_w0[188][3:0]) | ({4{loc_sram_buff_w1[188][4]}} & loc_sram_buff_w1[188][3:0]) | ({4{loc_sram_buff_w2[188][4]}} & loc_sram_buff_w2[188][3:0]) | ({4{loc_sram_buff_w3[188][4]}} & loc_sram_buff_w3[188][3:0]) | ({4{loc_sram_buff_w4[188][4]}} & loc_sram_buff_w4[188][3:0]) | ({4{loc_sram_buff_w5[188][4]}} & loc_sram_buff_w5[188][3:0]) | ({4{loc_sram_buff_w6[188][4]}} & loc_sram_buff_w6[188][3:0]) | ({4{loc_sram_buff_w7[188][4]}} & loc_sram_buff_w7[188][3:0]) | ({4{loc_sram_buff_w8[188][4]}} & loc_sram_buff_w8[188][3:0]) | ({4{loc_sram_buff_w9[188][4]}} & loc_sram_buff_w9[188][3:0]) | ({4{loc_sram_buff_w10[188][4]}} & loc_sram_buff_w10[188][3:0]) | ({4{loc_sram_buff_w11[188][4]}} & loc_sram_buff_w11[188][3:0]) | ({4{loc_sram_buff_w12[188][4]}} & loc_sram_buff_w12[188][3:0]) | ({4{loc_sram_buff_w13[188][4]}} & loc_sram_buff_w13[188][3:0]) | ({4{loc_sram_buff_w14[188][4]}} & loc_sram_buff_w14[188][3:0]) | ({4{loc_sram_buff_w15[188][4]}} & loc_sram_buff_w15[188][3:0]);
	loc_rdata_buff[ 267: 264] = ({4{loc_sram_buff_w0[189][4]}} & loc_sram_buff_w0[189][3:0]) | ({4{loc_sram_buff_w1[189][4]}} & loc_sram_buff_w1[189][3:0]) | ({4{loc_sram_buff_w2[189][4]}} & loc_sram_buff_w2[189][3:0]) | ({4{loc_sram_buff_w3[189][4]}} & loc_sram_buff_w3[189][3:0]) | ({4{loc_sram_buff_w4[189][4]}} & loc_sram_buff_w4[189][3:0]) | ({4{loc_sram_buff_w5[189][4]}} & loc_sram_buff_w5[189][3:0]) | ({4{loc_sram_buff_w6[189][4]}} & loc_sram_buff_w6[189][3:0]) | ({4{loc_sram_buff_w7[189][4]}} & loc_sram_buff_w7[189][3:0]) | ({4{loc_sram_buff_w8[189][4]}} & loc_sram_buff_w8[189][3:0]) | ({4{loc_sram_buff_w9[189][4]}} & loc_sram_buff_w9[189][3:0]) | ({4{loc_sram_buff_w10[189][4]}} & loc_sram_buff_w10[189][3:0]) | ({4{loc_sram_buff_w11[189][4]}} & loc_sram_buff_w11[189][3:0]) | ({4{loc_sram_buff_w12[189][4]}} & loc_sram_buff_w12[189][3:0]) | ({4{loc_sram_buff_w13[189][4]}} & loc_sram_buff_w13[189][3:0]) | ({4{loc_sram_buff_w14[189][4]}} & loc_sram_buff_w14[189][3:0]) | ({4{loc_sram_buff_w15[189][4]}} & loc_sram_buff_w15[189][3:0]);
	loc_rdata_buff[ 263: 260] = ({4{loc_sram_buff_w0[190][4]}} & loc_sram_buff_w0[190][3:0]) | ({4{loc_sram_buff_w1[190][4]}} & loc_sram_buff_w1[190][3:0]) | ({4{loc_sram_buff_w2[190][4]}} & loc_sram_buff_w2[190][3:0]) | ({4{loc_sram_buff_w3[190][4]}} & loc_sram_buff_w3[190][3:0]) | ({4{loc_sram_buff_w4[190][4]}} & loc_sram_buff_w4[190][3:0]) | ({4{loc_sram_buff_w5[190][4]}} & loc_sram_buff_w5[190][3:0]) | ({4{loc_sram_buff_w6[190][4]}} & loc_sram_buff_w6[190][3:0]) | ({4{loc_sram_buff_w7[190][4]}} & loc_sram_buff_w7[190][3:0]) | ({4{loc_sram_buff_w8[190][4]}} & loc_sram_buff_w8[190][3:0]) | ({4{loc_sram_buff_w9[190][4]}} & loc_sram_buff_w9[190][3:0]) | ({4{loc_sram_buff_w10[190][4]}} & loc_sram_buff_w10[190][3:0]) | ({4{loc_sram_buff_w11[190][4]}} & loc_sram_buff_w11[190][3:0]) | ({4{loc_sram_buff_w12[190][4]}} & loc_sram_buff_w12[190][3:0]) | ({4{loc_sram_buff_w13[190][4]}} & loc_sram_buff_w13[190][3:0]) | ({4{loc_sram_buff_w14[190][4]}} & loc_sram_buff_w14[190][3:0]) | ({4{loc_sram_buff_w15[190][4]}} & loc_sram_buff_w15[190][3:0]);
	loc_rdata_buff[ 259: 256] = ({4{loc_sram_buff_w0[191][4]}} & loc_sram_buff_w0[191][3:0]) | ({4{loc_sram_buff_w1[191][4]}} & loc_sram_buff_w1[191][3:0]) | ({4{loc_sram_buff_w2[191][4]}} & loc_sram_buff_w2[191][3:0]) | ({4{loc_sram_buff_w3[191][4]}} & loc_sram_buff_w3[191][3:0]) | ({4{loc_sram_buff_w4[191][4]}} & loc_sram_buff_w4[191][3:0]) | ({4{loc_sram_buff_w5[191][4]}} & loc_sram_buff_w5[191][3:0]) | ({4{loc_sram_buff_w6[191][4]}} & loc_sram_buff_w6[191][3:0]) | ({4{loc_sram_buff_w7[191][4]}} & loc_sram_buff_w7[191][3:0]) | ({4{loc_sram_buff_w8[191][4]}} & loc_sram_buff_w8[191][3:0]) | ({4{loc_sram_buff_w9[191][4]}} & loc_sram_buff_w9[191][3:0]) | ({4{loc_sram_buff_w10[191][4]}} & loc_sram_buff_w10[191][3:0]) | ({4{loc_sram_buff_w11[191][4]}} & loc_sram_buff_w11[191][3:0]) | ({4{loc_sram_buff_w12[191][4]}} & loc_sram_buff_w12[191][3:0]) | ({4{loc_sram_buff_w13[191][4]}} & loc_sram_buff_w13[191][3:0]) | ({4{loc_sram_buff_w14[191][4]}} & loc_sram_buff_w14[191][3:0]) | ({4{loc_sram_buff_w15[191][4]}} & loc_sram_buff_w15[191][3:0]);
	loc_rdata_buff[ 255: 252] = ({4{loc_sram_buff_w0[192][4]}} & loc_sram_buff_w0[192][3:0]) | ({4{loc_sram_buff_w1[192][4]}} & loc_sram_buff_w1[192][3:0]) | ({4{loc_sram_buff_w2[192][4]}} & loc_sram_buff_w2[192][3:0]) | ({4{loc_sram_buff_w3[192][4]}} & loc_sram_buff_w3[192][3:0]) | ({4{loc_sram_buff_w4[192][4]}} & loc_sram_buff_w4[192][3:0]) | ({4{loc_sram_buff_w5[192][4]}} & loc_sram_buff_w5[192][3:0]) | ({4{loc_sram_buff_w6[192][4]}} & loc_sram_buff_w6[192][3:0]) | ({4{loc_sram_buff_w7[192][4]}} & loc_sram_buff_w7[192][3:0]) | ({4{loc_sram_buff_w8[192][4]}} & loc_sram_buff_w8[192][3:0]) | ({4{loc_sram_buff_w9[192][4]}} & loc_sram_buff_w9[192][3:0]) | ({4{loc_sram_buff_w10[192][4]}} & loc_sram_buff_w10[192][3:0]) | ({4{loc_sram_buff_w11[192][4]}} & loc_sram_buff_w11[192][3:0]) | ({4{loc_sram_buff_w12[192][4]}} & loc_sram_buff_w12[192][3:0]) | ({4{loc_sram_buff_w13[192][4]}} & loc_sram_buff_w13[192][3:0]) | ({4{loc_sram_buff_w14[192][4]}} & loc_sram_buff_w14[192][3:0]) | ({4{loc_sram_buff_w15[192][4]}} & loc_sram_buff_w15[192][3:0]);
	loc_rdata_buff[ 251: 248] = ({4{loc_sram_buff_w0[193][4]}} & loc_sram_buff_w0[193][3:0]) | ({4{loc_sram_buff_w1[193][4]}} & loc_sram_buff_w1[193][3:0]) | ({4{loc_sram_buff_w2[193][4]}} & loc_sram_buff_w2[193][3:0]) | ({4{loc_sram_buff_w3[193][4]}} & loc_sram_buff_w3[193][3:0]) | ({4{loc_sram_buff_w4[193][4]}} & loc_sram_buff_w4[193][3:0]) | ({4{loc_sram_buff_w5[193][4]}} & loc_sram_buff_w5[193][3:0]) | ({4{loc_sram_buff_w6[193][4]}} & loc_sram_buff_w6[193][3:0]) | ({4{loc_sram_buff_w7[193][4]}} & loc_sram_buff_w7[193][3:0]) | ({4{loc_sram_buff_w8[193][4]}} & loc_sram_buff_w8[193][3:0]) | ({4{loc_sram_buff_w9[193][4]}} & loc_sram_buff_w9[193][3:0]) | ({4{loc_sram_buff_w10[193][4]}} & loc_sram_buff_w10[193][3:0]) | ({4{loc_sram_buff_w11[193][4]}} & loc_sram_buff_w11[193][3:0]) | ({4{loc_sram_buff_w12[193][4]}} & loc_sram_buff_w12[193][3:0]) | ({4{loc_sram_buff_w13[193][4]}} & loc_sram_buff_w13[193][3:0]) | ({4{loc_sram_buff_w14[193][4]}} & loc_sram_buff_w14[193][3:0]) | ({4{loc_sram_buff_w15[193][4]}} & loc_sram_buff_w15[193][3:0]);
	loc_rdata_buff[ 247: 244] = ({4{loc_sram_buff_w0[194][4]}} & loc_sram_buff_w0[194][3:0]) | ({4{loc_sram_buff_w1[194][4]}} & loc_sram_buff_w1[194][3:0]) | ({4{loc_sram_buff_w2[194][4]}} & loc_sram_buff_w2[194][3:0]) | ({4{loc_sram_buff_w3[194][4]}} & loc_sram_buff_w3[194][3:0]) | ({4{loc_sram_buff_w4[194][4]}} & loc_sram_buff_w4[194][3:0]) | ({4{loc_sram_buff_w5[194][4]}} & loc_sram_buff_w5[194][3:0]) | ({4{loc_sram_buff_w6[194][4]}} & loc_sram_buff_w6[194][3:0]) | ({4{loc_sram_buff_w7[194][4]}} & loc_sram_buff_w7[194][3:0]) | ({4{loc_sram_buff_w8[194][4]}} & loc_sram_buff_w8[194][3:0]) | ({4{loc_sram_buff_w9[194][4]}} & loc_sram_buff_w9[194][3:0]) | ({4{loc_sram_buff_w10[194][4]}} & loc_sram_buff_w10[194][3:0]) | ({4{loc_sram_buff_w11[194][4]}} & loc_sram_buff_w11[194][3:0]) | ({4{loc_sram_buff_w12[194][4]}} & loc_sram_buff_w12[194][3:0]) | ({4{loc_sram_buff_w13[194][4]}} & loc_sram_buff_w13[194][3:0]) | ({4{loc_sram_buff_w14[194][4]}} & loc_sram_buff_w14[194][3:0]) | ({4{loc_sram_buff_w15[194][4]}} & loc_sram_buff_w15[194][3:0]);
	loc_rdata_buff[ 243: 240] = ({4{loc_sram_buff_w0[195][4]}} & loc_sram_buff_w0[195][3:0]) | ({4{loc_sram_buff_w1[195][4]}} & loc_sram_buff_w1[195][3:0]) | ({4{loc_sram_buff_w2[195][4]}} & loc_sram_buff_w2[195][3:0]) | ({4{loc_sram_buff_w3[195][4]}} & loc_sram_buff_w3[195][3:0]) | ({4{loc_sram_buff_w4[195][4]}} & loc_sram_buff_w4[195][3:0]) | ({4{loc_sram_buff_w5[195][4]}} & loc_sram_buff_w5[195][3:0]) | ({4{loc_sram_buff_w6[195][4]}} & loc_sram_buff_w6[195][3:0]) | ({4{loc_sram_buff_w7[195][4]}} & loc_sram_buff_w7[195][3:0]) | ({4{loc_sram_buff_w8[195][4]}} & loc_sram_buff_w8[195][3:0]) | ({4{loc_sram_buff_w9[195][4]}} & loc_sram_buff_w9[195][3:0]) | ({4{loc_sram_buff_w10[195][4]}} & loc_sram_buff_w10[195][3:0]) | ({4{loc_sram_buff_w11[195][4]}} & loc_sram_buff_w11[195][3:0]) | ({4{loc_sram_buff_w12[195][4]}} & loc_sram_buff_w12[195][3:0]) | ({4{loc_sram_buff_w13[195][4]}} & loc_sram_buff_w13[195][3:0]) | ({4{loc_sram_buff_w14[195][4]}} & loc_sram_buff_w14[195][3:0]) | ({4{loc_sram_buff_w15[195][4]}} & loc_sram_buff_w15[195][3:0]);
	loc_rdata_buff[ 239: 236] = ({4{loc_sram_buff_w0[196][4]}} & loc_sram_buff_w0[196][3:0]) | ({4{loc_sram_buff_w1[196][4]}} & loc_sram_buff_w1[196][3:0]) | ({4{loc_sram_buff_w2[196][4]}} & loc_sram_buff_w2[196][3:0]) | ({4{loc_sram_buff_w3[196][4]}} & loc_sram_buff_w3[196][3:0]) | ({4{loc_sram_buff_w4[196][4]}} & loc_sram_buff_w4[196][3:0]) | ({4{loc_sram_buff_w5[196][4]}} & loc_sram_buff_w5[196][3:0]) | ({4{loc_sram_buff_w6[196][4]}} & loc_sram_buff_w6[196][3:0]) | ({4{loc_sram_buff_w7[196][4]}} & loc_sram_buff_w7[196][3:0]) | ({4{loc_sram_buff_w8[196][4]}} & loc_sram_buff_w8[196][3:0]) | ({4{loc_sram_buff_w9[196][4]}} & loc_sram_buff_w9[196][3:0]) | ({4{loc_sram_buff_w10[196][4]}} & loc_sram_buff_w10[196][3:0]) | ({4{loc_sram_buff_w11[196][4]}} & loc_sram_buff_w11[196][3:0]) | ({4{loc_sram_buff_w12[196][4]}} & loc_sram_buff_w12[196][3:0]) | ({4{loc_sram_buff_w13[196][4]}} & loc_sram_buff_w13[196][3:0]) | ({4{loc_sram_buff_w14[196][4]}} & loc_sram_buff_w14[196][3:0]) | ({4{loc_sram_buff_w15[196][4]}} & loc_sram_buff_w15[196][3:0]);
	loc_rdata_buff[ 235: 232] = ({4{loc_sram_buff_w0[197][4]}} & loc_sram_buff_w0[197][3:0]) | ({4{loc_sram_buff_w1[197][4]}} & loc_sram_buff_w1[197][3:0]) | ({4{loc_sram_buff_w2[197][4]}} & loc_sram_buff_w2[197][3:0]) | ({4{loc_sram_buff_w3[197][4]}} & loc_sram_buff_w3[197][3:0]) | ({4{loc_sram_buff_w4[197][4]}} & loc_sram_buff_w4[197][3:0]) | ({4{loc_sram_buff_w5[197][4]}} & loc_sram_buff_w5[197][3:0]) | ({4{loc_sram_buff_w6[197][4]}} & loc_sram_buff_w6[197][3:0]) | ({4{loc_sram_buff_w7[197][4]}} & loc_sram_buff_w7[197][3:0]) | ({4{loc_sram_buff_w8[197][4]}} & loc_sram_buff_w8[197][3:0]) | ({4{loc_sram_buff_w9[197][4]}} & loc_sram_buff_w9[197][3:0]) | ({4{loc_sram_buff_w10[197][4]}} & loc_sram_buff_w10[197][3:0]) | ({4{loc_sram_buff_w11[197][4]}} & loc_sram_buff_w11[197][3:0]) | ({4{loc_sram_buff_w12[197][4]}} & loc_sram_buff_w12[197][3:0]) | ({4{loc_sram_buff_w13[197][4]}} & loc_sram_buff_w13[197][3:0]) | ({4{loc_sram_buff_w14[197][4]}} & loc_sram_buff_w14[197][3:0]) | ({4{loc_sram_buff_w15[197][4]}} & loc_sram_buff_w15[197][3:0]);
	loc_rdata_buff[ 231: 228] = ({4{loc_sram_buff_w0[198][4]}} & loc_sram_buff_w0[198][3:0]) | ({4{loc_sram_buff_w1[198][4]}} & loc_sram_buff_w1[198][3:0]) | ({4{loc_sram_buff_w2[198][4]}} & loc_sram_buff_w2[198][3:0]) | ({4{loc_sram_buff_w3[198][4]}} & loc_sram_buff_w3[198][3:0]) | ({4{loc_sram_buff_w4[198][4]}} & loc_sram_buff_w4[198][3:0]) | ({4{loc_sram_buff_w5[198][4]}} & loc_sram_buff_w5[198][3:0]) | ({4{loc_sram_buff_w6[198][4]}} & loc_sram_buff_w6[198][3:0]) | ({4{loc_sram_buff_w7[198][4]}} & loc_sram_buff_w7[198][3:0]) | ({4{loc_sram_buff_w8[198][4]}} & loc_sram_buff_w8[198][3:0]) | ({4{loc_sram_buff_w9[198][4]}} & loc_sram_buff_w9[198][3:0]) | ({4{loc_sram_buff_w10[198][4]}} & loc_sram_buff_w10[198][3:0]) | ({4{loc_sram_buff_w11[198][4]}} & loc_sram_buff_w11[198][3:0]) | ({4{loc_sram_buff_w12[198][4]}} & loc_sram_buff_w12[198][3:0]) | ({4{loc_sram_buff_w13[198][4]}} & loc_sram_buff_w13[198][3:0]) | ({4{loc_sram_buff_w14[198][4]}} & loc_sram_buff_w14[198][3:0]) | ({4{loc_sram_buff_w15[198][4]}} & loc_sram_buff_w15[198][3:0]);
	loc_rdata_buff[ 227: 224] = ({4{loc_sram_buff_w0[199][4]}} & loc_sram_buff_w0[199][3:0]) | ({4{loc_sram_buff_w1[199][4]}} & loc_sram_buff_w1[199][3:0]) | ({4{loc_sram_buff_w2[199][4]}} & loc_sram_buff_w2[199][3:0]) | ({4{loc_sram_buff_w3[199][4]}} & loc_sram_buff_w3[199][3:0]) | ({4{loc_sram_buff_w4[199][4]}} & loc_sram_buff_w4[199][3:0]) | ({4{loc_sram_buff_w5[199][4]}} & loc_sram_buff_w5[199][3:0]) | ({4{loc_sram_buff_w6[199][4]}} & loc_sram_buff_w6[199][3:0]) | ({4{loc_sram_buff_w7[199][4]}} & loc_sram_buff_w7[199][3:0]) | ({4{loc_sram_buff_w8[199][4]}} & loc_sram_buff_w8[199][3:0]) | ({4{loc_sram_buff_w9[199][4]}} & loc_sram_buff_w9[199][3:0]) | ({4{loc_sram_buff_w10[199][4]}} & loc_sram_buff_w10[199][3:0]) | ({4{loc_sram_buff_w11[199][4]}} & loc_sram_buff_w11[199][3:0]) | ({4{loc_sram_buff_w12[199][4]}} & loc_sram_buff_w12[199][3:0]) | ({4{loc_sram_buff_w13[199][4]}} & loc_sram_buff_w13[199][3:0]) | ({4{loc_sram_buff_w14[199][4]}} & loc_sram_buff_w14[199][3:0]) | ({4{loc_sram_buff_w15[199][4]}} & loc_sram_buff_w15[199][3:0]);
	loc_rdata_buff[ 223: 220] = ({4{loc_sram_buff_w0[200][4]}} & loc_sram_buff_w0[200][3:0]) | ({4{loc_sram_buff_w1[200][4]}} & loc_sram_buff_w1[200][3:0]) | ({4{loc_sram_buff_w2[200][4]}} & loc_sram_buff_w2[200][3:0]) | ({4{loc_sram_buff_w3[200][4]}} & loc_sram_buff_w3[200][3:0]) | ({4{loc_sram_buff_w4[200][4]}} & loc_sram_buff_w4[200][3:0]) | ({4{loc_sram_buff_w5[200][4]}} & loc_sram_buff_w5[200][3:0]) | ({4{loc_sram_buff_w6[200][4]}} & loc_sram_buff_w6[200][3:0]) | ({4{loc_sram_buff_w7[200][4]}} & loc_sram_buff_w7[200][3:0]) | ({4{loc_sram_buff_w8[200][4]}} & loc_sram_buff_w8[200][3:0]) | ({4{loc_sram_buff_w9[200][4]}} & loc_sram_buff_w9[200][3:0]) | ({4{loc_sram_buff_w10[200][4]}} & loc_sram_buff_w10[200][3:0]) | ({4{loc_sram_buff_w11[200][4]}} & loc_sram_buff_w11[200][3:0]) | ({4{loc_sram_buff_w12[200][4]}} & loc_sram_buff_w12[200][3:0]) | ({4{loc_sram_buff_w13[200][4]}} & loc_sram_buff_w13[200][3:0]) | ({4{loc_sram_buff_w14[200][4]}} & loc_sram_buff_w14[200][3:0]) | ({4{loc_sram_buff_w15[200][4]}} & loc_sram_buff_w15[200][3:0]);
	loc_rdata_buff[ 219: 216] = ({4{loc_sram_buff_w0[201][4]}} & loc_sram_buff_w0[201][3:0]) | ({4{loc_sram_buff_w1[201][4]}} & loc_sram_buff_w1[201][3:0]) | ({4{loc_sram_buff_w2[201][4]}} & loc_sram_buff_w2[201][3:0]) | ({4{loc_sram_buff_w3[201][4]}} & loc_sram_buff_w3[201][3:0]) | ({4{loc_sram_buff_w4[201][4]}} & loc_sram_buff_w4[201][3:0]) | ({4{loc_sram_buff_w5[201][4]}} & loc_sram_buff_w5[201][3:0]) | ({4{loc_sram_buff_w6[201][4]}} & loc_sram_buff_w6[201][3:0]) | ({4{loc_sram_buff_w7[201][4]}} & loc_sram_buff_w7[201][3:0]) | ({4{loc_sram_buff_w8[201][4]}} & loc_sram_buff_w8[201][3:0]) | ({4{loc_sram_buff_w9[201][4]}} & loc_sram_buff_w9[201][3:0]) | ({4{loc_sram_buff_w10[201][4]}} & loc_sram_buff_w10[201][3:0]) | ({4{loc_sram_buff_w11[201][4]}} & loc_sram_buff_w11[201][3:0]) | ({4{loc_sram_buff_w12[201][4]}} & loc_sram_buff_w12[201][3:0]) | ({4{loc_sram_buff_w13[201][4]}} & loc_sram_buff_w13[201][3:0]) | ({4{loc_sram_buff_w14[201][4]}} & loc_sram_buff_w14[201][3:0]) | ({4{loc_sram_buff_w15[201][4]}} & loc_sram_buff_w15[201][3:0]);
	loc_rdata_buff[ 215: 212] = ({4{loc_sram_buff_w0[202][4]}} & loc_sram_buff_w0[202][3:0]) | ({4{loc_sram_buff_w1[202][4]}} & loc_sram_buff_w1[202][3:0]) | ({4{loc_sram_buff_w2[202][4]}} & loc_sram_buff_w2[202][3:0]) | ({4{loc_sram_buff_w3[202][4]}} & loc_sram_buff_w3[202][3:0]) | ({4{loc_sram_buff_w4[202][4]}} & loc_sram_buff_w4[202][3:0]) | ({4{loc_sram_buff_w5[202][4]}} & loc_sram_buff_w5[202][3:0]) | ({4{loc_sram_buff_w6[202][4]}} & loc_sram_buff_w6[202][3:0]) | ({4{loc_sram_buff_w7[202][4]}} & loc_sram_buff_w7[202][3:0]) | ({4{loc_sram_buff_w8[202][4]}} & loc_sram_buff_w8[202][3:0]) | ({4{loc_sram_buff_w9[202][4]}} & loc_sram_buff_w9[202][3:0]) | ({4{loc_sram_buff_w10[202][4]}} & loc_sram_buff_w10[202][3:0]) | ({4{loc_sram_buff_w11[202][4]}} & loc_sram_buff_w11[202][3:0]) | ({4{loc_sram_buff_w12[202][4]}} & loc_sram_buff_w12[202][3:0]) | ({4{loc_sram_buff_w13[202][4]}} & loc_sram_buff_w13[202][3:0]) | ({4{loc_sram_buff_w14[202][4]}} & loc_sram_buff_w14[202][3:0]) | ({4{loc_sram_buff_w15[202][4]}} & loc_sram_buff_w15[202][3:0]);
	loc_rdata_buff[ 211: 208] = ({4{loc_sram_buff_w0[203][4]}} & loc_sram_buff_w0[203][3:0]) | ({4{loc_sram_buff_w1[203][4]}} & loc_sram_buff_w1[203][3:0]) | ({4{loc_sram_buff_w2[203][4]}} & loc_sram_buff_w2[203][3:0]) | ({4{loc_sram_buff_w3[203][4]}} & loc_sram_buff_w3[203][3:0]) | ({4{loc_sram_buff_w4[203][4]}} & loc_sram_buff_w4[203][3:0]) | ({4{loc_sram_buff_w5[203][4]}} & loc_sram_buff_w5[203][3:0]) | ({4{loc_sram_buff_w6[203][4]}} & loc_sram_buff_w6[203][3:0]) | ({4{loc_sram_buff_w7[203][4]}} & loc_sram_buff_w7[203][3:0]) | ({4{loc_sram_buff_w8[203][4]}} & loc_sram_buff_w8[203][3:0]) | ({4{loc_sram_buff_w9[203][4]}} & loc_sram_buff_w9[203][3:0]) | ({4{loc_sram_buff_w10[203][4]}} & loc_sram_buff_w10[203][3:0]) | ({4{loc_sram_buff_w11[203][4]}} & loc_sram_buff_w11[203][3:0]) | ({4{loc_sram_buff_w12[203][4]}} & loc_sram_buff_w12[203][3:0]) | ({4{loc_sram_buff_w13[203][4]}} & loc_sram_buff_w13[203][3:0]) | ({4{loc_sram_buff_w14[203][4]}} & loc_sram_buff_w14[203][3:0]) | ({4{loc_sram_buff_w15[203][4]}} & loc_sram_buff_w15[203][3:0]);
	loc_rdata_buff[ 207: 204] = ({4{loc_sram_buff_w0[204][4]}} & loc_sram_buff_w0[204][3:0]) | ({4{loc_sram_buff_w1[204][4]}} & loc_sram_buff_w1[204][3:0]) | ({4{loc_sram_buff_w2[204][4]}} & loc_sram_buff_w2[204][3:0]) | ({4{loc_sram_buff_w3[204][4]}} & loc_sram_buff_w3[204][3:0]) | ({4{loc_sram_buff_w4[204][4]}} & loc_sram_buff_w4[204][3:0]) | ({4{loc_sram_buff_w5[204][4]}} & loc_sram_buff_w5[204][3:0]) | ({4{loc_sram_buff_w6[204][4]}} & loc_sram_buff_w6[204][3:0]) | ({4{loc_sram_buff_w7[204][4]}} & loc_sram_buff_w7[204][3:0]) | ({4{loc_sram_buff_w8[204][4]}} & loc_sram_buff_w8[204][3:0]) | ({4{loc_sram_buff_w9[204][4]}} & loc_sram_buff_w9[204][3:0]) | ({4{loc_sram_buff_w10[204][4]}} & loc_sram_buff_w10[204][3:0]) | ({4{loc_sram_buff_w11[204][4]}} & loc_sram_buff_w11[204][3:0]) | ({4{loc_sram_buff_w12[204][4]}} & loc_sram_buff_w12[204][3:0]) | ({4{loc_sram_buff_w13[204][4]}} & loc_sram_buff_w13[204][3:0]) | ({4{loc_sram_buff_w14[204][4]}} & loc_sram_buff_w14[204][3:0]) | ({4{loc_sram_buff_w15[204][4]}} & loc_sram_buff_w15[204][3:0]);
	loc_rdata_buff[ 203: 200] = ({4{loc_sram_buff_w0[205][4]}} & loc_sram_buff_w0[205][3:0]) | ({4{loc_sram_buff_w1[205][4]}} & loc_sram_buff_w1[205][3:0]) | ({4{loc_sram_buff_w2[205][4]}} & loc_sram_buff_w2[205][3:0]) | ({4{loc_sram_buff_w3[205][4]}} & loc_sram_buff_w3[205][3:0]) | ({4{loc_sram_buff_w4[205][4]}} & loc_sram_buff_w4[205][3:0]) | ({4{loc_sram_buff_w5[205][4]}} & loc_sram_buff_w5[205][3:0]) | ({4{loc_sram_buff_w6[205][4]}} & loc_sram_buff_w6[205][3:0]) | ({4{loc_sram_buff_w7[205][4]}} & loc_sram_buff_w7[205][3:0]) | ({4{loc_sram_buff_w8[205][4]}} & loc_sram_buff_w8[205][3:0]) | ({4{loc_sram_buff_w9[205][4]}} & loc_sram_buff_w9[205][3:0]) | ({4{loc_sram_buff_w10[205][4]}} & loc_sram_buff_w10[205][3:0]) | ({4{loc_sram_buff_w11[205][4]}} & loc_sram_buff_w11[205][3:0]) | ({4{loc_sram_buff_w12[205][4]}} & loc_sram_buff_w12[205][3:0]) | ({4{loc_sram_buff_w13[205][4]}} & loc_sram_buff_w13[205][3:0]) | ({4{loc_sram_buff_w14[205][4]}} & loc_sram_buff_w14[205][3:0]) | ({4{loc_sram_buff_w15[205][4]}} & loc_sram_buff_w15[205][3:0]);
	loc_rdata_buff[ 199: 196] = ({4{loc_sram_buff_w0[206][4]}} & loc_sram_buff_w0[206][3:0]) | ({4{loc_sram_buff_w1[206][4]}} & loc_sram_buff_w1[206][3:0]) | ({4{loc_sram_buff_w2[206][4]}} & loc_sram_buff_w2[206][3:0]) | ({4{loc_sram_buff_w3[206][4]}} & loc_sram_buff_w3[206][3:0]) | ({4{loc_sram_buff_w4[206][4]}} & loc_sram_buff_w4[206][3:0]) | ({4{loc_sram_buff_w5[206][4]}} & loc_sram_buff_w5[206][3:0]) | ({4{loc_sram_buff_w6[206][4]}} & loc_sram_buff_w6[206][3:0]) | ({4{loc_sram_buff_w7[206][4]}} & loc_sram_buff_w7[206][3:0]) | ({4{loc_sram_buff_w8[206][4]}} & loc_sram_buff_w8[206][3:0]) | ({4{loc_sram_buff_w9[206][4]}} & loc_sram_buff_w9[206][3:0]) | ({4{loc_sram_buff_w10[206][4]}} & loc_sram_buff_w10[206][3:0]) | ({4{loc_sram_buff_w11[206][4]}} & loc_sram_buff_w11[206][3:0]) | ({4{loc_sram_buff_w12[206][4]}} & loc_sram_buff_w12[206][3:0]) | ({4{loc_sram_buff_w13[206][4]}} & loc_sram_buff_w13[206][3:0]) | ({4{loc_sram_buff_w14[206][4]}} & loc_sram_buff_w14[206][3:0]) | ({4{loc_sram_buff_w15[206][4]}} & loc_sram_buff_w15[206][3:0]);
	loc_rdata_buff[ 195: 192] = ({4{loc_sram_buff_w0[207][4]}} & loc_sram_buff_w0[207][3:0]) | ({4{loc_sram_buff_w1[207][4]}} & loc_sram_buff_w1[207][3:0]) | ({4{loc_sram_buff_w2[207][4]}} & loc_sram_buff_w2[207][3:0]) | ({4{loc_sram_buff_w3[207][4]}} & loc_sram_buff_w3[207][3:0]) | ({4{loc_sram_buff_w4[207][4]}} & loc_sram_buff_w4[207][3:0]) | ({4{loc_sram_buff_w5[207][4]}} & loc_sram_buff_w5[207][3:0]) | ({4{loc_sram_buff_w6[207][4]}} & loc_sram_buff_w6[207][3:0]) | ({4{loc_sram_buff_w7[207][4]}} & loc_sram_buff_w7[207][3:0]) | ({4{loc_sram_buff_w8[207][4]}} & loc_sram_buff_w8[207][3:0]) | ({4{loc_sram_buff_w9[207][4]}} & loc_sram_buff_w9[207][3:0]) | ({4{loc_sram_buff_w10[207][4]}} & loc_sram_buff_w10[207][3:0]) | ({4{loc_sram_buff_w11[207][4]}} & loc_sram_buff_w11[207][3:0]) | ({4{loc_sram_buff_w12[207][4]}} & loc_sram_buff_w12[207][3:0]) | ({4{loc_sram_buff_w13[207][4]}} & loc_sram_buff_w13[207][3:0]) | ({4{loc_sram_buff_w14[207][4]}} & loc_sram_buff_w14[207][3:0]) | ({4{loc_sram_buff_w15[207][4]}} & loc_sram_buff_w15[207][3:0]);
	loc_rdata_buff[ 191: 188] = ({4{loc_sram_buff_w0[208][4]}} & loc_sram_buff_w0[208][3:0]) | ({4{loc_sram_buff_w1[208][4]}} & loc_sram_buff_w1[208][3:0]) | ({4{loc_sram_buff_w2[208][4]}} & loc_sram_buff_w2[208][3:0]) | ({4{loc_sram_buff_w3[208][4]}} & loc_sram_buff_w3[208][3:0]) | ({4{loc_sram_buff_w4[208][4]}} & loc_sram_buff_w4[208][3:0]) | ({4{loc_sram_buff_w5[208][4]}} & loc_sram_buff_w5[208][3:0]) | ({4{loc_sram_buff_w6[208][4]}} & loc_sram_buff_w6[208][3:0]) | ({4{loc_sram_buff_w7[208][4]}} & loc_sram_buff_w7[208][3:0]) | ({4{loc_sram_buff_w8[208][4]}} & loc_sram_buff_w8[208][3:0]) | ({4{loc_sram_buff_w9[208][4]}} & loc_sram_buff_w9[208][3:0]) | ({4{loc_sram_buff_w10[208][4]}} & loc_sram_buff_w10[208][3:0]) | ({4{loc_sram_buff_w11[208][4]}} & loc_sram_buff_w11[208][3:0]) | ({4{loc_sram_buff_w12[208][4]}} & loc_sram_buff_w12[208][3:0]) | ({4{loc_sram_buff_w13[208][4]}} & loc_sram_buff_w13[208][3:0]) | ({4{loc_sram_buff_w14[208][4]}} & loc_sram_buff_w14[208][3:0]) | ({4{loc_sram_buff_w15[208][4]}} & loc_sram_buff_w15[208][3:0]);
	loc_rdata_buff[ 187: 184] = ({4{loc_sram_buff_w0[209][4]}} & loc_sram_buff_w0[209][3:0]) | ({4{loc_sram_buff_w1[209][4]}} & loc_sram_buff_w1[209][3:0]) | ({4{loc_sram_buff_w2[209][4]}} & loc_sram_buff_w2[209][3:0]) | ({4{loc_sram_buff_w3[209][4]}} & loc_sram_buff_w3[209][3:0]) | ({4{loc_sram_buff_w4[209][4]}} & loc_sram_buff_w4[209][3:0]) | ({4{loc_sram_buff_w5[209][4]}} & loc_sram_buff_w5[209][3:0]) | ({4{loc_sram_buff_w6[209][4]}} & loc_sram_buff_w6[209][3:0]) | ({4{loc_sram_buff_w7[209][4]}} & loc_sram_buff_w7[209][3:0]) | ({4{loc_sram_buff_w8[209][4]}} & loc_sram_buff_w8[209][3:0]) | ({4{loc_sram_buff_w9[209][4]}} & loc_sram_buff_w9[209][3:0]) | ({4{loc_sram_buff_w10[209][4]}} & loc_sram_buff_w10[209][3:0]) | ({4{loc_sram_buff_w11[209][4]}} & loc_sram_buff_w11[209][3:0]) | ({4{loc_sram_buff_w12[209][4]}} & loc_sram_buff_w12[209][3:0]) | ({4{loc_sram_buff_w13[209][4]}} & loc_sram_buff_w13[209][3:0]) | ({4{loc_sram_buff_w14[209][4]}} & loc_sram_buff_w14[209][3:0]) | ({4{loc_sram_buff_w15[209][4]}} & loc_sram_buff_w15[209][3:0]);
	loc_rdata_buff[ 183: 180] = ({4{loc_sram_buff_w0[210][4]}} & loc_sram_buff_w0[210][3:0]) | ({4{loc_sram_buff_w1[210][4]}} & loc_sram_buff_w1[210][3:0]) | ({4{loc_sram_buff_w2[210][4]}} & loc_sram_buff_w2[210][3:0]) | ({4{loc_sram_buff_w3[210][4]}} & loc_sram_buff_w3[210][3:0]) | ({4{loc_sram_buff_w4[210][4]}} & loc_sram_buff_w4[210][3:0]) | ({4{loc_sram_buff_w5[210][4]}} & loc_sram_buff_w5[210][3:0]) | ({4{loc_sram_buff_w6[210][4]}} & loc_sram_buff_w6[210][3:0]) | ({4{loc_sram_buff_w7[210][4]}} & loc_sram_buff_w7[210][3:0]) | ({4{loc_sram_buff_w8[210][4]}} & loc_sram_buff_w8[210][3:0]) | ({4{loc_sram_buff_w9[210][4]}} & loc_sram_buff_w9[210][3:0]) | ({4{loc_sram_buff_w10[210][4]}} & loc_sram_buff_w10[210][3:0]) | ({4{loc_sram_buff_w11[210][4]}} & loc_sram_buff_w11[210][3:0]) | ({4{loc_sram_buff_w12[210][4]}} & loc_sram_buff_w12[210][3:0]) | ({4{loc_sram_buff_w13[210][4]}} & loc_sram_buff_w13[210][3:0]) | ({4{loc_sram_buff_w14[210][4]}} & loc_sram_buff_w14[210][3:0]) | ({4{loc_sram_buff_w15[210][4]}} & loc_sram_buff_w15[210][3:0]);
	loc_rdata_buff[ 179: 176] = ({4{loc_sram_buff_w0[211][4]}} & loc_sram_buff_w0[211][3:0]) | ({4{loc_sram_buff_w1[211][4]}} & loc_sram_buff_w1[211][3:0]) | ({4{loc_sram_buff_w2[211][4]}} & loc_sram_buff_w2[211][3:0]) | ({4{loc_sram_buff_w3[211][4]}} & loc_sram_buff_w3[211][3:0]) | ({4{loc_sram_buff_w4[211][4]}} & loc_sram_buff_w4[211][3:0]) | ({4{loc_sram_buff_w5[211][4]}} & loc_sram_buff_w5[211][3:0]) | ({4{loc_sram_buff_w6[211][4]}} & loc_sram_buff_w6[211][3:0]) | ({4{loc_sram_buff_w7[211][4]}} & loc_sram_buff_w7[211][3:0]) | ({4{loc_sram_buff_w8[211][4]}} & loc_sram_buff_w8[211][3:0]) | ({4{loc_sram_buff_w9[211][4]}} & loc_sram_buff_w9[211][3:0]) | ({4{loc_sram_buff_w10[211][4]}} & loc_sram_buff_w10[211][3:0]) | ({4{loc_sram_buff_w11[211][4]}} & loc_sram_buff_w11[211][3:0]) | ({4{loc_sram_buff_w12[211][4]}} & loc_sram_buff_w12[211][3:0]) | ({4{loc_sram_buff_w13[211][4]}} & loc_sram_buff_w13[211][3:0]) | ({4{loc_sram_buff_w14[211][4]}} & loc_sram_buff_w14[211][3:0]) | ({4{loc_sram_buff_w15[211][4]}} & loc_sram_buff_w15[211][3:0]);
	loc_rdata_buff[ 175: 172] = ({4{loc_sram_buff_w0[212][4]}} & loc_sram_buff_w0[212][3:0]) | ({4{loc_sram_buff_w1[212][4]}} & loc_sram_buff_w1[212][3:0]) | ({4{loc_sram_buff_w2[212][4]}} & loc_sram_buff_w2[212][3:0]) | ({4{loc_sram_buff_w3[212][4]}} & loc_sram_buff_w3[212][3:0]) | ({4{loc_sram_buff_w4[212][4]}} & loc_sram_buff_w4[212][3:0]) | ({4{loc_sram_buff_w5[212][4]}} & loc_sram_buff_w5[212][3:0]) | ({4{loc_sram_buff_w6[212][4]}} & loc_sram_buff_w6[212][3:0]) | ({4{loc_sram_buff_w7[212][4]}} & loc_sram_buff_w7[212][3:0]) | ({4{loc_sram_buff_w8[212][4]}} & loc_sram_buff_w8[212][3:0]) | ({4{loc_sram_buff_w9[212][4]}} & loc_sram_buff_w9[212][3:0]) | ({4{loc_sram_buff_w10[212][4]}} & loc_sram_buff_w10[212][3:0]) | ({4{loc_sram_buff_w11[212][4]}} & loc_sram_buff_w11[212][3:0]) | ({4{loc_sram_buff_w12[212][4]}} & loc_sram_buff_w12[212][3:0]) | ({4{loc_sram_buff_w13[212][4]}} & loc_sram_buff_w13[212][3:0]) | ({4{loc_sram_buff_w14[212][4]}} & loc_sram_buff_w14[212][3:0]) | ({4{loc_sram_buff_w15[212][4]}} & loc_sram_buff_w15[212][3:0]);
	loc_rdata_buff[ 171: 168] = ({4{loc_sram_buff_w0[213][4]}} & loc_sram_buff_w0[213][3:0]) | ({4{loc_sram_buff_w1[213][4]}} & loc_sram_buff_w1[213][3:0]) | ({4{loc_sram_buff_w2[213][4]}} & loc_sram_buff_w2[213][3:0]) | ({4{loc_sram_buff_w3[213][4]}} & loc_sram_buff_w3[213][3:0]) | ({4{loc_sram_buff_w4[213][4]}} & loc_sram_buff_w4[213][3:0]) | ({4{loc_sram_buff_w5[213][4]}} & loc_sram_buff_w5[213][3:0]) | ({4{loc_sram_buff_w6[213][4]}} & loc_sram_buff_w6[213][3:0]) | ({4{loc_sram_buff_w7[213][4]}} & loc_sram_buff_w7[213][3:0]) | ({4{loc_sram_buff_w8[213][4]}} & loc_sram_buff_w8[213][3:0]) | ({4{loc_sram_buff_w9[213][4]}} & loc_sram_buff_w9[213][3:0]) | ({4{loc_sram_buff_w10[213][4]}} & loc_sram_buff_w10[213][3:0]) | ({4{loc_sram_buff_w11[213][4]}} & loc_sram_buff_w11[213][3:0]) | ({4{loc_sram_buff_w12[213][4]}} & loc_sram_buff_w12[213][3:0]) | ({4{loc_sram_buff_w13[213][4]}} & loc_sram_buff_w13[213][3:0]) | ({4{loc_sram_buff_w14[213][4]}} & loc_sram_buff_w14[213][3:0]) | ({4{loc_sram_buff_w15[213][4]}} & loc_sram_buff_w15[213][3:0]);
	loc_rdata_buff[ 167: 164] = ({4{loc_sram_buff_w0[214][4]}} & loc_sram_buff_w0[214][3:0]) | ({4{loc_sram_buff_w1[214][4]}} & loc_sram_buff_w1[214][3:0]) | ({4{loc_sram_buff_w2[214][4]}} & loc_sram_buff_w2[214][3:0]) | ({4{loc_sram_buff_w3[214][4]}} & loc_sram_buff_w3[214][3:0]) | ({4{loc_sram_buff_w4[214][4]}} & loc_sram_buff_w4[214][3:0]) | ({4{loc_sram_buff_w5[214][4]}} & loc_sram_buff_w5[214][3:0]) | ({4{loc_sram_buff_w6[214][4]}} & loc_sram_buff_w6[214][3:0]) | ({4{loc_sram_buff_w7[214][4]}} & loc_sram_buff_w7[214][3:0]) | ({4{loc_sram_buff_w8[214][4]}} & loc_sram_buff_w8[214][3:0]) | ({4{loc_sram_buff_w9[214][4]}} & loc_sram_buff_w9[214][3:0]) | ({4{loc_sram_buff_w10[214][4]}} & loc_sram_buff_w10[214][3:0]) | ({4{loc_sram_buff_w11[214][4]}} & loc_sram_buff_w11[214][3:0]) | ({4{loc_sram_buff_w12[214][4]}} & loc_sram_buff_w12[214][3:0]) | ({4{loc_sram_buff_w13[214][4]}} & loc_sram_buff_w13[214][3:0]) | ({4{loc_sram_buff_w14[214][4]}} & loc_sram_buff_w14[214][3:0]) | ({4{loc_sram_buff_w15[214][4]}} & loc_sram_buff_w15[214][3:0]);
	loc_rdata_buff[ 163: 160] = ({4{loc_sram_buff_w0[215][4]}} & loc_sram_buff_w0[215][3:0]) | ({4{loc_sram_buff_w1[215][4]}} & loc_sram_buff_w1[215][3:0]) | ({4{loc_sram_buff_w2[215][4]}} & loc_sram_buff_w2[215][3:0]) | ({4{loc_sram_buff_w3[215][4]}} & loc_sram_buff_w3[215][3:0]) | ({4{loc_sram_buff_w4[215][4]}} & loc_sram_buff_w4[215][3:0]) | ({4{loc_sram_buff_w5[215][4]}} & loc_sram_buff_w5[215][3:0]) | ({4{loc_sram_buff_w6[215][4]}} & loc_sram_buff_w6[215][3:0]) | ({4{loc_sram_buff_w7[215][4]}} & loc_sram_buff_w7[215][3:0]) | ({4{loc_sram_buff_w8[215][4]}} & loc_sram_buff_w8[215][3:0]) | ({4{loc_sram_buff_w9[215][4]}} & loc_sram_buff_w9[215][3:0]) | ({4{loc_sram_buff_w10[215][4]}} & loc_sram_buff_w10[215][3:0]) | ({4{loc_sram_buff_w11[215][4]}} & loc_sram_buff_w11[215][3:0]) | ({4{loc_sram_buff_w12[215][4]}} & loc_sram_buff_w12[215][3:0]) | ({4{loc_sram_buff_w13[215][4]}} & loc_sram_buff_w13[215][3:0]) | ({4{loc_sram_buff_w14[215][4]}} & loc_sram_buff_w14[215][3:0]) | ({4{loc_sram_buff_w15[215][4]}} & loc_sram_buff_w15[215][3:0]);
	loc_rdata_buff[ 159: 156] = ({4{loc_sram_buff_w0[216][4]}} & loc_sram_buff_w0[216][3:0]) | ({4{loc_sram_buff_w1[216][4]}} & loc_sram_buff_w1[216][3:0]) | ({4{loc_sram_buff_w2[216][4]}} & loc_sram_buff_w2[216][3:0]) | ({4{loc_sram_buff_w3[216][4]}} & loc_sram_buff_w3[216][3:0]) | ({4{loc_sram_buff_w4[216][4]}} & loc_sram_buff_w4[216][3:0]) | ({4{loc_sram_buff_w5[216][4]}} & loc_sram_buff_w5[216][3:0]) | ({4{loc_sram_buff_w6[216][4]}} & loc_sram_buff_w6[216][3:0]) | ({4{loc_sram_buff_w7[216][4]}} & loc_sram_buff_w7[216][3:0]) | ({4{loc_sram_buff_w8[216][4]}} & loc_sram_buff_w8[216][3:0]) | ({4{loc_sram_buff_w9[216][4]}} & loc_sram_buff_w9[216][3:0]) | ({4{loc_sram_buff_w10[216][4]}} & loc_sram_buff_w10[216][3:0]) | ({4{loc_sram_buff_w11[216][4]}} & loc_sram_buff_w11[216][3:0]) | ({4{loc_sram_buff_w12[216][4]}} & loc_sram_buff_w12[216][3:0]) | ({4{loc_sram_buff_w13[216][4]}} & loc_sram_buff_w13[216][3:0]) | ({4{loc_sram_buff_w14[216][4]}} & loc_sram_buff_w14[216][3:0]) | ({4{loc_sram_buff_w15[216][4]}} & loc_sram_buff_w15[216][3:0]);
	loc_rdata_buff[ 155: 152] = ({4{loc_sram_buff_w0[217][4]}} & loc_sram_buff_w0[217][3:0]) | ({4{loc_sram_buff_w1[217][4]}} & loc_sram_buff_w1[217][3:0]) | ({4{loc_sram_buff_w2[217][4]}} & loc_sram_buff_w2[217][3:0]) | ({4{loc_sram_buff_w3[217][4]}} & loc_sram_buff_w3[217][3:0]) | ({4{loc_sram_buff_w4[217][4]}} & loc_sram_buff_w4[217][3:0]) | ({4{loc_sram_buff_w5[217][4]}} & loc_sram_buff_w5[217][3:0]) | ({4{loc_sram_buff_w6[217][4]}} & loc_sram_buff_w6[217][3:0]) | ({4{loc_sram_buff_w7[217][4]}} & loc_sram_buff_w7[217][3:0]) | ({4{loc_sram_buff_w8[217][4]}} & loc_sram_buff_w8[217][3:0]) | ({4{loc_sram_buff_w9[217][4]}} & loc_sram_buff_w9[217][3:0]) | ({4{loc_sram_buff_w10[217][4]}} & loc_sram_buff_w10[217][3:0]) | ({4{loc_sram_buff_w11[217][4]}} & loc_sram_buff_w11[217][3:0]) | ({4{loc_sram_buff_w12[217][4]}} & loc_sram_buff_w12[217][3:0]) | ({4{loc_sram_buff_w13[217][4]}} & loc_sram_buff_w13[217][3:0]) | ({4{loc_sram_buff_w14[217][4]}} & loc_sram_buff_w14[217][3:0]) | ({4{loc_sram_buff_w15[217][4]}} & loc_sram_buff_w15[217][3:0]);
	loc_rdata_buff[ 151: 148] = ({4{loc_sram_buff_w0[218][4]}} & loc_sram_buff_w0[218][3:0]) | ({4{loc_sram_buff_w1[218][4]}} & loc_sram_buff_w1[218][3:0]) | ({4{loc_sram_buff_w2[218][4]}} & loc_sram_buff_w2[218][3:0]) | ({4{loc_sram_buff_w3[218][4]}} & loc_sram_buff_w3[218][3:0]) | ({4{loc_sram_buff_w4[218][4]}} & loc_sram_buff_w4[218][3:0]) | ({4{loc_sram_buff_w5[218][4]}} & loc_sram_buff_w5[218][3:0]) | ({4{loc_sram_buff_w6[218][4]}} & loc_sram_buff_w6[218][3:0]) | ({4{loc_sram_buff_w7[218][4]}} & loc_sram_buff_w7[218][3:0]) | ({4{loc_sram_buff_w8[218][4]}} & loc_sram_buff_w8[218][3:0]) | ({4{loc_sram_buff_w9[218][4]}} & loc_sram_buff_w9[218][3:0]) | ({4{loc_sram_buff_w10[218][4]}} & loc_sram_buff_w10[218][3:0]) | ({4{loc_sram_buff_w11[218][4]}} & loc_sram_buff_w11[218][3:0]) | ({4{loc_sram_buff_w12[218][4]}} & loc_sram_buff_w12[218][3:0]) | ({4{loc_sram_buff_w13[218][4]}} & loc_sram_buff_w13[218][3:0]) | ({4{loc_sram_buff_w14[218][4]}} & loc_sram_buff_w14[218][3:0]) | ({4{loc_sram_buff_w15[218][4]}} & loc_sram_buff_w15[218][3:0]);
	loc_rdata_buff[ 147: 144] = ({4{loc_sram_buff_w0[219][4]}} & loc_sram_buff_w0[219][3:0]) | ({4{loc_sram_buff_w1[219][4]}} & loc_sram_buff_w1[219][3:0]) | ({4{loc_sram_buff_w2[219][4]}} & loc_sram_buff_w2[219][3:0]) | ({4{loc_sram_buff_w3[219][4]}} & loc_sram_buff_w3[219][3:0]) | ({4{loc_sram_buff_w4[219][4]}} & loc_sram_buff_w4[219][3:0]) | ({4{loc_sram_buff_w5[219][4]}} & loc_sram_buff_w5[219][3:0]) | ({4{loc_sram_buff_w6[219][4]}} & loc_sram_buff_w6[219][3:0]) | ({4{loc_sram_buff_w7[219][4]}} & loc_sram_buff_w7[219][3:0]) | ({4{loc_sram_buff_w8[219][4]}} & loc_sram_buff_w8[219][3:0]) | ({4{loc_sram_buff_w9[219][4]}} & loc_sram_buff_w9[219][3:0]) | ({4{loc_sram_buff_w10[219][4]}} & loc_sram_buff_w10[219][3:0]) | ({4{loc_sram_buff_w11[219][4]}} & loc_sram_buff_w11[219][3:0]) | ({4{loc_sram_buff_w12[219][4]}} & loc_sram_buff_w12[219][3:0]) | ({4{loc_sram_buff_w13[219][4]}} & loc_sram_buff_w13[219][3:0]) | ({4{loc_sram_buff_w14[219][4]}} & loc_sram_buff_w14[219][3:0]) | ({4{loc_sram_buff_w15[219][4]}} & loc_sram_buff_w15[219][3:0]);
	loc_rdata_buff[ 143: 140] = ({4{loc_sram_buff_w0[220][4]}} & loc_sram_buff_w0[220][3:0]) | ({4{loc_sram_buff_w1[220][4]}} & loc_sram_buff_w1[220][3:0]) | ({4{loc_sram_buff_w2[220][4]}} & loc_sram_buff_w2[220][3:0]) | ({4{loc_sram_buff_w3[220][4]}} & loc_sram_buff_w3[220][3:0]) | ({4{loc_sram_buff_w4[220][4]}} & loc_sram_buff_w4[220][3:0]) | ({4{loc_sram_buff_w5[220][4]}} & loc_sram_buff_w5[220][3:0]) | ({4{loc_sram_buff_w6[220][4]}} & loc_sram_buff_w6[220][3:0]) | ({4{loc_sram_buff_w7[220][4]}} & loc_sram_buff_w7[220][3:0]) | ({4{loc_sram_buff_w8[220][4]}} & loc_sram_buff_w8[220][3:0]) | ({4{loc_sram_buff_w9[220][4]}} & loc_sram_buff_w9[220][3:0]) | ({4{loc_sram_buff_w10[220][4]}} & loc_sram_buff_w10[220][3:0]) | ({4{loc_sram_buff_w11[220][4]}} & loc_sram_buff_w11[220][3:0]) | ({4{loc_sram_buff_w12[220][4]}} & loc_sram_buff_w12[220][3:0]) | ({4{loc_sram_buff_w13[220][4]}} & loc_sram_buff_w13[220][3:0]) | ({4{loc_sram_buff_w14[220][4]}} & loc_sram_buff_w14[220][3:0]) | ({4{loc_sram_buff_w15[220][4]}} & loc_sram_buff_w15[220][3:0]);
	loc_rdata_buff[ 139: 136] = ({4{loc_sram_buff_w0[221][4]}} & loc_sram_buff_w0[221][3:0]) | ({4{loc_sram_buff_w1[221][4]}} & loc_sram_buff_w1[221][3:0]) | ({4{loc_sram_buff_w2[221][4]}} & loc_sram_buff_w2[221][3:0]) | ({4{loc_sram_buff_w3[221][4]}} & loc_sram_buff_w3[221][3:0]) | ({4{loc_sram_buff_w4[221][4]}} & loc_sram_buff_w4[221][3:0]) | ({4{loc_sram_buff_w5[221][4]}} & loc_sram_buff_w5[221][3:0]) | ({4{loc_sram_buff_w6[221][4]}} & loc_sram_buff_w6[221][3:0]) | ({4{loc_sram_buff_w7[221][4]}} & loc_sram_buff_w7[221][3:0]) | ({4{loc_sram_buff_w8[221][4]}} & loc_sram_buff_w8[221][3:0]) | ({4{loc_sram_buff_w9[221][4]}} & loc_sram_buff_w9[221][3:0]) | ({4{loc_sram_buff_w10[221][4]}} & loc_sram_buff_w10[221][3:0]) | ({4{loc_sram_buff_w11[221][4]}} & loc_sram_buff_w11[221][3:0]) | ({4{loc_sram_buff_w12[221][4]}} & loc_sram_buff_w12[221][3:0]) | ({4{loc_sram_buff_w13[221][4]}} & loc_sram_buff_w13[221][3:0]) | ({4{loc_sram_buff_w14[221][4]}} & loc_sram_buff_w14[221][3:0]) | ({4{loc_sram_buff_w15[221][4]}} & loc_sram_buff_w15[221][3:0]);
	loc_rdata_buff[ 135: 132] = ({4{loc_sram_buff_w0[222][4]}} & loc_sram_buff_w0[222][3:0]) | ({4{loc_sram_buff_w1[222][4]}} & loc_sram_buff_w1[222][3:0]) | ({4{loc_sram_buff_w2[222][4]}} & loc_sram_buff_w2[222][3:0]) | ({4{loc_sram_buff_w3[222][4]}} & loc_sram_buff_w3[222][3:0]) | ({4{loc_sram_buff_w4[222][4]}} & loc_sram_buff_w4[222][3:0]) | ({4{loc_sram_buff_w5[222][4]}} & loc_sram_buff_w5[222][3:0]) | ({4{loc_sram_buff_w6[222][4]}} & loc_sram_buff_w6[222][3:0]) | ({4{loc_sram_buff_w7[222][4]}} & loc_sram_buff_w7[222][3:0]) | ({4{loc_sram_buff_w8[222][4]}} & loc_sram_buff_w8[222][3:0]) | ({4{loc_sram_buff_w9[222][4]}} & loc_sram_buff_w9[222][3:0]) | ({4{loc_sram_buff_w10[222][4]}} & loc_sram_buff_w10[222][3:0]) | ({4{loc_sram_buff_w11[222][4]}} & loc_sram_buff_w11[222][3:0]) | ({4{loc_sram_buff_w12[222][4]}} & loc_sram_buff_w12[222][3:0]) | ({4{loc_sram_buff_w13[222][4]}} & loc_sram_buff_w13[222][3:0]) | ({4{loc_sram_buff_w14[222][4]}} & loc_sram_buff_w14[222][3:0]) | ({4{loc_sram_buff_w15[222][4]}} & loc_sram_buff_w15[222][3:0]);
	loc_rdata_buff[ 131: 128] = ({4{loc_sram_buff_w0[223][4]}} & loc_sram_buff_w0[223][3:0]) | ({4{loc_sram_buff_w1[223][4]}} & loc_sram_buff_w1[223][3:0]) | ({4{loc_sram_buff_w2[223][4]}} & loc_sram_buff_w2[223][3:0]) | ({4{loc_sram_buff_w3[223][4]}} & loc_sram_buff_w3[223][3:0]) | ({4{loc_sram_buff_w4[223][4]}} & loc_sram_buff_w4[223][3:0]) | ({4{loc_sram_buff_w5[223][4]}} & loc_sram_buff_w5[223][3:0]) | ({4{loc_sram_buff_w6[223][4]}} & loc_sram_buff_w6[223][3:0]) | ({4{loc_sram_buff_w7[223][4]}} & loc_sram_buff_w7[223][3:0]) | ({4{loc_sram_buff_w8[223][4]}} & loc_sram_buff_w8[223][3:0]) | ({4{loc_sram_buff_w9[223][4]}} & loc_sram_buff_w9[223][3:0]) | ({4{loc_sram_buff_w10[223][4]}} & loc_sram_buff_w10[223][3:0]) | ({4{loc_sram_buff_w11[223][4]}} & loc_sram_buff_w11[223][3:0]) | ({4{loc_sram_buff_w12[223][4]}} & loc_sram_buff_w12[223][3:0]) | ({4{loc_sram_buff_w13[223][4]}} & loc_sram_buff_w13[223][3:0]) | ({4{loc_sram_buff_w14[223][4]}} & loc_sram_buff_w14[223][3:0]) | ({4{loc_sram_buff_w15[223][4]}} & loc_sram_buff_w15[223][3:0]);
	loc_rdata_buff[ 127: 124] = ({4{loc_sram_buff_w0[224][4]}} & loc_sram_buff_w0[224][3:0]) | ({4{loc_sram_buff_w1[224][4]}} & loc_sram_buff_w1[224][3:0]) | ({4{loc_sram_buff_w2[224][4]}} & loc_sram_buff_w2[224][3:0]) | ({4{loc_sram_buff_w3[224][4]}} & loc_sram_buff_w3[224][3:0]) | ({4{loc_sram_buff_w4[224][4]}} & loc_sram_buff_w4[224][3:0]) | ({4{loc_sram_buff_w5[224][4]}} & loc_sram_buff_w5[224][3:0]) | ({4{loc_sram_buff_w6[224][4]}} & loc_sram_buff_w6[224][3:0]) | ({4{loc_sram_buff_w7[224][4]}} & loc_sram_buff_w7[224][3:0]) | ({4{loc_sram_buff_w8[224][4]}} & loc_sram_buff_w8[224][3:0]) | ({4{loc_sram_buff_w9[224][4]}} & loc_sram_buff_w9[224][3:0]) | ({4{loc_sram_buff_w10[224][4]}} & loc_sram_buff_w10[224][3:0]) | ({4{loc_sram_buff_w11[224][4]}} & loc_sram_buff_w11[224][3:0]) | ({4{loc_sram_buff_w12[224][4]}} & loc_sram_buff_w12[224][3:0]) | ({4{loc_sram_buff_w13[224][4]}} & loc_sram_buff_w13[224][3:0]) | ({4{loc_sram_buff_w14[224][4]}} & loc_sram_buff_w14[224][3:0]) | ({4{loc_sram_buff_w15[224][4]}} & loc_sram_buff_w15[224][3:0]);
	loc_rdata_buff[ 123: 120] = ({4{loc_sram_buff_w0[225][4]}} & loc_sram_buff_w0[225][3:0]) | ({4{loc_sram_buff_w1[225][4]}} & loc_sram_buff_w1[225][3:0]) | ({4{loc_sram_buff_w2[225][4]}} & loc_sram_buff_w2[225][3:0]) | ({4{loc_sram_buff_w3[225][4]}} & loc_sram_buff_w3[225][3:0]) | ({4{loc_sram_buff_w4[225][4]}} & loc_sram_buff_w4[225][3:0]) | ({4{loc_sram_buff_w5[225][4]}} & loc_sram_buff_w5[225][3:0]) | ({4{loc_sram_buff_w6[225][4]}} & loc_sram_buff_w6[225][3:0]) | ({4{loc_sram_buff_w7[225][4]}} & loc_sram_buff_w7[225][3:0]) | ({4{loc_sram_buff_w8[225][4]}} & loc_sram_buff_w8[225][3:0]) | ({4{loc_sram_buff_w9[225][4]}} & loc_sram_buff_w9[225][3:0]) | ({4{loc_sram_buff_w10[225][4]}} & loc_sram_buff_w10[225][3:0]) | ({4{loc_sram_buff_w11[225][4]}} & loc_sram_buff_w11[225][3:0]) | ({4{loc_sram_buff_w12[225][4]}} & loc_sram_buff_w12[225][3:0]) | ({4{loc_sram_buff_w13[225][4]}} & loc_sram_buff_w13[225][3:0]) | ({4{loc_sram_buff_w14[225][4]}} & loc_sram_buff_w14[225][3:0]) | ({4{loc_sram_buff_w15[225][4]}} & loc_sram_buff_w15[225][3:0]);
	loc_rdata_buff[ 119: 116] = ({4{loc_sram_buff_w0[226][4]}} & loc_sram_buff_w0[226][3:0]) | ({4{loc_sram_buff_w1[226][4]}} & loc_sram_buff_w1[226][3:0]) | ({4{loc_sram_buff_w2[226][4]}} & loc_sram_buff_w2[226][3:0]) | ({4{loc_sram_buff_w3[226][4]}} & loc_sram_buff_w3[226][3:0]) | ({4{loc_sram_buff_w4[226][4]}} & loc_sram_buff_w4[226][3:0]) | ({4{loc_sram_buff_w5[226][4]}} & loc_sram_buff_w5[226][3:0]) | ({4{loc_sram_buff_w6[226][4]}} & loc_sram_buff_w6[226][3:0]) | ({4{loc_sram_buff_w7[226][4]}} & loc_sram_buff_w7[226][3:0]) | ({4{loc_sram_buff_w8[226][4]}} & loc_sram_buff_w8[226][3:0]) | ({4{loc_sram_buff_w9[226][4]}} & loc_sram_buff_w9[226][3:0]) | ({4{loc_sram_buff_w10[226][4]}} & loc_sram_buff_w10[226][3:0]) | ({4{loc_sram_buff_w11[226][4]}} & loc_sram_buff_w11[226][3:0]) | ({4{loc_sram_buff_w12[226][4]}} & loc_sram_buff_w12[226][3:0]) | ({4{loc_sram_buff_w13[226][4]}} & loc_sram_buff_w13[226][3:0]) | ({4{loc_sram_buff_w14[226][4]}} & loc_sram_buff_w14[226][3:0]) | ({4{loc_sram_buff_w15[226][4]}} & loc_sram_buff_w15[226][3:0]);
	loc_rdata_buff[ 115: 112] = ({4{loc_sram_buff_w0[227][4]}} & loc_sram_buff_w0[227][3:0]) | ({4{loc_sram_buff_w1[227][4]}} & loc_sram_buff_w1[227][3:0]) | ({4{loc_sram_buff_w2[227][4]}} & loc_sram_buff_w2[227][3:0]) | ({4{loc_sram_buff_w3[227][4]}} & loc_sram_buff_w3[227][3:0]) | ({4{loc_sram_buff_w4[227][4]}} & loc_sram_buff_w4[227][3:0]) | ({4{loc_sram_buff_w5[227][4]}} & loc_sram_buff_w5[227][3:0]) | ({4{loc_sram_buff_w6[227][4]}} & loc_sram_buff_w6[227][3:0]) | ({4{loc_sram_buff_w7[227][4]}} & loc_sram_buff_w7[227][3:0]) | ({4{loc_sram_buff_w8[227][4]}} & loc_sram_buff_w8[227][3:0]) | ({4{loc_sram_buff_w9[227][4]}} & loc_sram_buff_w9[227][3:0]) | ({4{loc_sram_buff_w10[227][4]}} & loc_sram_buff_w10[227][3:0]) | ({4{loc_sram_buff_w11[227][4]}} & loc_sram_buff_w11[227][3:0]) | ({4{loc_sram_buff_w12[227][4]}} & loc_sram_buff_w12[227][3:0]) | ({4{loc_sram_buff_w13[227][4]}} & loc_sram_buff_w13[227][3:0]) | ({4{loc_sram_buff_w14[227][4]}} & loc_sram_buff_w14[227][3:0]) | ({4{loc_sram_buff_w15[227][4]}} & loc_sram_buff_w15[227][3:0]);
	loc_rdata_buff[ 111: 108] = ({4{loc_sram_buff_w0[228][4]}} & loc_sram_buff_w0[228][3:0]) | ({4{loc_sram_buff_w1[228][4]}} & loc_sram_buff_w1[228][3:0]) | ({4{loc_sram_buff_w2[228][4]}} & loc_sram_buff_w2[228][3:0]) | ({4{loc_sram_buff_w3[228][4]}} & loc_sram_buff_w3[228][3:0]) | ({4{loc_sram_buff_w4[228][4]}} & loc_sram_buff_w4[228][3:0]) | ({4{loc_sram_buff_w5[228][4]}} & loc_sram_buff_w5[228][3:0]) | ({4{loc_sram_buff_w6[228][4]}} & loc_sram_buff_w6[228][3:0]) | ({4{loc_sram_buff_w7[228][4]}} & loc_sram_buff_w7[228][3:0]) | ({4{loc_sram_buff_w8[228][4]}} & loc_sram_buff_w8[228][3:0]) | ({4{loc_sram_buff_w9[228][4]}} & loc_sram_buff_w9[228][3:0]) | ({4{loc_sram_buff_w10[228][4]}} & loc_sram_buff_w10[228][3:0]) | ({4{loc_sram_buff_w11[228][4]}} & loc_sram_buff_w11[228][3:0]) | ({4{loc_sram_buff_w12[228][4]}} & loc_sram_buff_w12[228][3:0]) | ({4{loc_sram_buff_w13[228][4]}} & loc_sram_buff_w13[228][3:0]) | ({4{loc_sram_buff_w14[228][4]}} & loc_sram_buff_w14[228][3:0]) | ({4{loc_sram_buff_w15[228][4]}} & loc_sram_buff_w15[228][3:0]);
	loc_rdata_buff[ 107: 104] = ({4{loc_sram_buff_w0[229][4]}} & loc_sram_buff_w0[229][3:0]) | ({4{loc_sram_buff_w1[229][4]}} & loc_sram_buff_w1[229][3:0]) | ({4{loc_sram_buff_w2[229][4]}} & loc_sram_buff_w2[229][3:0]) | ({4{loc_sram_buff_w3[229][4]}} & loc_sram_buff_w3[229][3:0]) | ({4{loc_sram_buff_w4[229][4]}} & loc_sram_buff_w4[229][3:0]) | ({4{loc_sram_buff_w5[229][4]}} & loc_sram_buff_w5[229][3:0]) | ({4{loc_sram_buff_w6[229][4]}} & loc_sram_buff_w6[229][3:0]) | ({4{loc_sram_buff_w7[229][4]}} & loc_sram_buff_w7[229][3:0]) | ({4{loc_sram_buff_w8[229][4]}} & loc_sram_buff_w8[229][3:0]) | ({4{loc_sram_buff_w9[229][4]}} & loc_sram_buff_w9[229][3:0]) | ({4{loc_sram_buff_w10[229][4]}} & loc_sram_buff_w10[229][3:0]) | ({4{loc_sram_buff_w11[229][4]}} & loc_sram_buff_w11[229][3:0]) | ({4{loc_sram_buff_w12[229][4]}} & loc_sram_buff_w12[229][3:0]) | ({4{loc_sram_buff_w13[229][4]}} & loc_sram_buff_w13[229][3:0]) | ({4{loc_sram_buff_w14[229][4]}} & loc_sram_buff_w14[229][3:0]) | ({4{loc_sram_buff_w15[229][4]}} & loc_sram_buff_w15[229][3:0]);
	loc_rdata_buff[ 103: 100] = ({4{loc_sram_buff_w0[230][4]}} & loc_sram_buff_w0[230][3:0]) | ({4{loc_sram_buff_w1[230][4]}} & loc_sram_buff_w1[230][3:0]) | ({4{loc_sram_buff_w2[230][4]}} & loc_sram_buff_w2[230][3:0]) | ({4{loc_sram_buff_w3[230][4]}} & loc_sram_buff_w3[230][3:0]) | ({4{loc_sram_buff_w4[230][4]}} & loc_sram_buff_w4[230][3:0]) | ({4{loc_sram_buff_w5[230][4]}} & loc_sram_buff_w5[230][3:0]) | ({4{loc_sram_buff_w6[230][4]}} & loc_sram_buff_w6[230][3:0]) | ({4{loc_sram_buff_w7[230][4]}} & loc_sram_buff_w7[230][3:0]) | ({4{loc_sram_buff_w8[230][4]}} & loc_sram_buff_w8[230][3:0]) | ({4{loc_sram_buff_w9[230][4]}} & loc_sram_buff_w9[230][3:0]) | ({4{loc_sram_buff_w10[230][4]}} & loc_sram_buff_w10[230][3:0]) | ({4{loc_sram_buff_w11[230][4]}} & loc_sram_buff_w11[230][3:0]) | ({4{loc_sram_buff_w12[230][4]}} & loc_sram_buff_w12[230][3:0]) | ({4{loc_sram_buff_w13[230][4]}} & loc_sram_buff_w13[230][3:0]) | ({4{loc_sram_buff_w14[230][4]}} & loc_sram_buff_w14[230][3:0]) | ({4{loc_sram_buff_w15[230][4]}} & loc_sram_buff_w15[230][3:0]);
	loc_rdata_buff[  99:  96] = ({4{loc_sram_buff_w0[231][4]}} & loc_sram_buff_w0[231][3:0]) | ({4{loc_sram_buff_w1[231][4]}} & loc_sram_buff_w1[231][3:0]) | ({4{loc_sram_buff_w2[231][4]}} & loc_sram_buff_w2[231][3:0]) | ({4{loc_sram_buff_w3[231][4]}} & loc_sram_buff_w3[231][3:0]) | ({4{loc_sram_buff_w4[231][4]}} & loc_sram_buff_w4[231][3:0]) | ({4{loc_sram_buff_w5[231][4]}} & loc_sram_buff_w5[231][3:0]) | ({4{loc_sram_buff_w6[231][4]}} & loc_sram_buff_w6[231][3:0]) | ({4{loc_sram_buff_w7[231][4]}} & loc_sram_buff_w7[231][3:0]) | ({4{loc_sram_buff_w8[231][4]}} & loc_sram_buff_w8[231][3:0]) | ({4{loc_sram_buff_w9[231][4]}} & loc_sram_buff_w9[231][3:0]) | ({4{loc_sram_buff_w10[231][4]}} & loc_sram_buff_w10[231][3:0]) | ({4{loc_sram_buff_w11[231][4]}} & loc_sram_buff_w11[231][3:0]) | ({4{loc_sram_buff_w12[231][4]}} & loc_sram_buff_w12[231][3:0]) | ({4{loc_sram_buff_w13[231][4]}} & loc_sram_buff_w13[231][3:0]) | ({4{loc_sram_buff_w14[231][4]}} & loc_sram_buff_w14[231][3:0]) | ({4{loc_sram_buff_w15[231][4]}} & loc_sram_buff_w15[231][3:0]);
	loc_rdata_buff[  95:  92] = ({4{loc_sram_buff_w0[232][4]}} & loc_sram_buff_w0[232][3:0]) | ({4{loc_sram_buff_w1[232][4]}} & loc_sram_buff_w1[232][3:0]) | ({4{loc_sram_buff_w2[232][4]}} & loc_sram_buff_w2[232][3:0]) | ({4{loc_sram_buff_w3[232][4]}} & loc_sram_buff_w3[232][3:0]) | ({4{loc_sram_buff_w4[232][4]}} & loc_sram_buff_w4[232][3:0]) | ({4{loc_sram_buff_w5[232][4]}} & loc_sram_buff_w5[232][3:0]) | ({4{loc_sram_buff_w6[232][4]}} & loc_sram_buff_w6[232][3:0]) | ({4{loc_sram_buff_w7[232][4]}} & loc_sram_buff_w7[232][3:0]) | ({4{loc_sram_buff_w8[232][4]}} & loc_sram_buff_w8[232][3:0]) | ({4{loc_sram_buff_w9[232][4]}} & loc_sram_buff_w9[232][3:0]) | ({4{loc_sram_buff_w10[232][4]}} & loc_sram_buff_w10[232][3:0]) | ({4{loc_sram_buff_w11[232][4]}} & loc_sram_buff_w11[232][3:0]) | ({4{loc_sram_buff_w12[232][4]}} & loc_sram_buff_w12[232][3:0]) | ({4{loc_sram_buff_w13[232][4]}} & loc_sram_buff_w13[232][3:0]) | ({4{loc_sram_buff_w14[232][4]}} & loc_sram_buff_w14[232][3:0]) | ({4{loc_sram_buff_w15[232][4]}} & loc_sram_buff_w15[232][3:0]);
	loc_rdata_buff[  91:  88] = ({4{loc_sram_buff_w0[233][4]}} & loc_sram_buff_w0[233][3:0]) | ({4{loc_sram_buff_w1[233][4]}} & loc_sram_buff_w1[233][3:0]) | ({4{loc_sram_buff_w2[233][4]}} & loc_sram_buff_w2[233][3:0]) | ({4{loc_sram_buff_w3[233][4]}} & loc_sram_buff_w3[233][3:0]) | ({4{loc_sram_buff_w4[233][4]}} & loc_sram_buff_w4[233][3:0]) | ({4{loc_sram_buff_w5[233][4]}} & loc_sram_buff_w5[233][3:0]) | ({4{loc_sram_buff_w6[233][4]}} & loc_sram_buff_w6[233][3:0]) | ({4{loc_sram_buff_w7[233][4]}} & loc_sram_buff_w7[233][3:0]) | ({4{loc_sram_buff_w8[233][4]}} & loc_sram_buff_w8[233][3:0]) | ({4{loc_sram_buff_w9[233][4]}} & loc_sram_buff_w9[233][3:0]) | ({4{loc_sram_buff_w10[233][4]}} & loc_sram_buff_w10[233][3:0]) | ({4{loc_sram_buff_w11[233][4]}} & loc_sram_buff_w11[233][3:0]) | ({4{loc_sram_buff_w12[233][4]}} & loc_sram_buff_w12[233][3:0]) | ({4{loc_sram_buff_w13[233][4]}} & loc_sram_buff_w13[233][3:0]) | ({4{loc_sram_buff_w14[233][4]}} & loc_sram_buff_w14[233][3:0]) | ({4{loc_sram_buff_w15[233][4]}} & loc_sram_buff_w15[233][3:0]);
	loc_rdata_buff[  87:  84] = ({4{loc_sram_buff_w0[234][4]}} & loc_sram_buff_w0[234][3:0]) | ({4{loc_sram_buff_w1[234][4]}} & loc_sram_buff_w1[234][3:0]) | ({4{loc_sram_buff_w2[234][4]}} & loc_sram_buff_w2[234][3:0]) | ({4{loc_sram_buff_w3[234][4]}} & loc_sram_buff_w3[234][3:0]) | ({4{loc_sram_buff_w4[234][4]}} & loc_sram_buff_w4[234][3:0]) | ({4{loc_sram_buff_w5[234][4]}} & loc_sram_buff_w5[234][3:0]) | ({4{loc_sram_buff_w6[234][4]}} & loc_sram_buff_w6[234][3:0]) | ({4{loc_sram_buff_w7[234][4]}} & loc_sram_buff_w7[234][3:0]) | ({4{loc_sram_buff_w8[234][4]}} & loc_sram_buff_w8[234][3:0]) | ({4{loc_sram_buff_w9[234][4]}} & loc_sram_buff_w9[234][3:0]) | ({4{loc_sram_buff_w10[234][4]}} & loc_sram_buff_w10[234][3:0]) | ({4{loc_sram_buff_w11[234][4]}} & loc_sram_buff_w11[234][3:0]) | ({4{loc_sram_buff_w12[234][4]}} & loc_sram_buff_w12[234][3:0]) | ({4{loc_sram_buff_w13[234][4]}} & loc_sram_buff_w13[234][3:0]) | ({4{loc_sram_buff_w14[234][4]}} & loc_sram_buff_w14[234][3:0]) | ({4{loc_sram_buff_w15[234][4]}} & loc_sram_buff_w15[234][3:0]);
	loc_rdata_buff[  83:  80] = ({4{loc_sram_buff_w0[235][4]}} & loc_sram_buff_w0[235][3:0]) | ({4{loc_sram_buff_w1[235][4]}} & loc_sram_buff_w1[235][3:0]) | ({4{loc_sram_buff_w2[235][4]}} & loc_sram_buff_w2[235][3:0]) | ({4{loc_sram_buff_w3[235][4]}} & loc_sram_buff_w3[235][3:0]) | ({4{loc_sram_buff_w4[235][4]}} & loc_sram_buff_w4[235][3:0]) | ({4{loc_sram_buff_w5[235][4]}} & loc_sram_buff_w5[235][3:0]) | ({4{loc_sram_buff_w6[235][4]}} & loc_sram_buff_w6[235][3:0]) | ({4{loc_sram_buff_w7[235][4]}} & loc_sram_buff_w7[235][3:0]) | ({4{loc_sram_buff_w8[235][4]}} & loc_sram_buff_w8[235][3:0]) | ({4{loc_sram_buff_w9[235][4]}} & loc_sram_buff_w9[235][3:0]) | ({4{loc_sram_buff_w10[235][4]}} & loc_sram_buff_w10[235][3:0]) | ({4{loc_sram_buff_w11[235][4]}} & loc_sram_buff_w11[235][3:0]) | ({4{loc_sram_buff_w12[235][4]}} & loc_sram_buff_w12[235][3:0]) | ({4{loc_sram_buff_w13[235][4]}} & loc_sram_buff_w13[235][3:0]) | ({4{loc_sram_buff_w14[235][4]}} & loc_sram_buff_w14[235][3:0]) | ({4{loc_sram_buff_w15[235][4]}} & loc_sram_buff_w15[235][3:0]);
	loc_rdata_buff[  79:  76] = ({4{loc_sram_buff_w0[236][4]}} & loc_sram_buff_w0[236][3:0]) | ({4{loc_sram_buff_w1[236][4]}} & loc_sram_buff_w1[236][3:0]) | ({4{loc_sram_buff_w2[236][4]}} & loc_sram_buff_w2[236][3:0]) | ({4{loc_sram_buff_w3[236][4]}} & loc_sram_buff_w3[236][3:0]) | ({4{loc_sram_buff_w4[236][4]}} & loc_sram_buff_w4[236][3:0]) | ({4{loc_sram_buff_w5[236][4]}} & loc_sram_buff_w5[236][3:0]) | ({4{loc_sram_buff_w6[236][4]}} & loc_sram_buff_w6[236][3:0]) | ({4{loc_sram_buff_w7[236][4]}} & loc_sram_buff_w7[236][3:0]) | ({4{loc_sram_buff_w8[236][4]}} & loc_sram_buff_w8[236][3:0]) | ({4{loc_sram_buff_w9[236][4]}} & loc_sram_buff_w9[236][3:0]) | ({4{loc_sram_buff_w10[236][4]}} & loc_sram_buff_w10[236][3:0]) | ({4{loc_sram_buff_w11[236][4]}} & loc_sram_buff_w11[236][3:0]) | ({4{loc_sram_buff_w12[236][4]}} & loc_sram_buff_w12[236][3:0]) | ({4{loc_sram_buff_w13[236][4]}} & loc_sram_buff_w13[236][3:0]) | ({4{loc_sram_buff_w14[236][4]}} & loc_sram_buff_w14[236][3:0]) | ({4{loc_sram_buff_w15[236][4]}} & loc_sram_buff_w15[236][3:0]);
	loc_rdata_buff[  75:  72] = ({4{loc_sram_buff_w0[237][4]}} & loc_sram_buff_w0[237][3:0]) | ({4{loc_sram_buff_w1[237][4]}} & loc_sram_buff_w1[237][3:0]) | ({4{loc_sram_buff_w2[237][4]}} & loc_sram_buff_w2[237][3:0]) | ({4{loc_sram_buff_w3[237][4]}} & loc_sram_buff_w3[237][3:0]) | ({4{loc_sram_buff_w4[237][4]}} & loc_sram_buff_w4[237][3:0]) | ({4{loc_sram_buff_w5[237][4]}} & loc_sram_buff_w5[237][3:0]) | ({4{loc_sram_buff_w6[237][4]}} & loc_sram_buff_w6[237][3:0]) | ({4{loc_sram_buff_w7[237][4]}} & loc_sram_buff_w7[237][3:0]) | ({4{loc_sram_buff_w8[237][4]}} & loc_sram_buff_w8[237][3:0]) | ({4{loc_sram_buff_w9[237][4]}} & loc_sram_buff_w9[237][3:0]) | ({4{loc_sram_buff_w10[237][4]}} & loc_sram_buff_w10[237][3:0]) | ({4{loc_sram_buff_w11[237][4]}} & loc_sram_buff_w11[237][3:0]) | ({4{loc_sram_buff_w12[237][4]}} & loc_sram_buff_w12[237][3:0]) | ({4{loc_sram_buff_w13[237][4]}} & loc_sram_buff_w13[237][3:0]) | ({4{loc_sram_buff_w14[237][4]}} & loc_sram_buff_w14[237][3:0]) | ({4{loc_sram_buff_w15[237][4]}} & loc_sram_buff_w15[237][3:0]);
	loc_rdata_buff[  71:  68] = ({4{loc_sram_buff_w0[238][4]}} & loc_sram_buff_w0[238][3:0]) | ({4{loc_sram_buff_w1[238][4]}} & loc_sram_buff_w1[238][3:0]) | ({4{loc_sram_buff_w2[238][4]}} & loc_sram_buff_w2[238][3:0]) | ({4{loc_sram_buff_w3[238][4]}} & loc_sram_buff_w3[238][3:0]) | ({4{loc_sram_buff_w4[238][4]}} & loc_sram_buff_w4[238][3:0]) | ({4{loc_sram_buff_w5[238][4]}} & loc_sram_buff_w5[238][3:0]) | ({4{loc_sram_buff_w6[238][4]}} & loc_sram_buff_w6[238][3:0]) | ({4{loc_sram_buff_w7[238][4]}} & loc_sram_buff_w7[238][3:0]) | ({4{loc_sram_buff_w8[238][4]}} & loc_sram_buff_w8[238][3:0]) | ({4{loc_sram_buff_w9[238][4]}} & loc_sram_buff_w9[238][3:0]) | ({4{loc_sram_buff_w10[238][4]}} & loc_sram_buff_w10[238][3:0]) | ({4{loc_sram_buff_w11[238][4]}} & loc_sram_buff_w11[238][3:0]) | ({4{loc_sram_buff_w12[238][4]}} & loc_sram_buff_w12[238][3:0]) | ({4{loc_sram_buff_w13[238][4]}} & loc_sram_buff_w13[238][3:0]) | ({4{loc_sram_buff_w14[238][4]}} & loc_sram_buff_w14[238][3:0]) | ({4{loc_sram_buff_w15[238][4]}} & loc_sram_buff_w15[238][3:0]);
	loc_rdata_buff[  67:  64] = ({4{loc_sram_buff_w0[239][4]}} & loc_sram_buff_w0[239][3:0]) | ({4{loc_sram_buff_w1[239][4]}} & loc_sram_buff_w1[239][3:0]) | ({4{loc_sram_buff_w2[239][4]}} & loc_sram_buff_w2[239][3:0]) | ({4{loc_sram_buff_w3[239][4]}} & loc_sram_buff_w3[239][3:0]) | ({4{loc_sram_buff_w4[239][4]}} & loc_sram_buff_w4[239][3:0]) | ({4{loc_sram_buff_w5[239][4]}} & loc_sram_buff_w5[239][3:0]) | ({4{loc_sram_buff_w6[239][4]}} & loc_sram_buff_w6[239][3:0]) | ({4{loc_sram_buff_w7[239][4]}} & loc_sram_buff_w7[239][3:0]) | ({4{loc_sram_buff_w8[239][4]}} & loc_sram_buff_w8[239][3:0]) | ({4{loc_sram_buff_w9[239][4]}} & loc_sram_buff_w9[239][3:0]) | ({4{loc_sram_buff_w10[239][4]}} & loc_sram_buff_w10[239][3:0]) | ({4{loc_sram_buff_w11[239][4]}} & loc_sram_buff_w11[239][3:0]) | ({4{loc_sram_buff_w12[239][4]}} & loc_sram_buff_w12[239][3:0]) | ({4{loc_sram_buff_w13[239][4]}} & loc_sram_buff_w13[239][3:0]) | ({4{loc_sram_buff_w14[239][4]}} & loc_sram_buff_w14[239][3:0]) | ({4{loc_sram_buff_w15[239][4]}} & loc_sram_buff_w15[239][3:0]);
	loc_rdata_buff[  63:  60] = ({4{loc_sram_buff_w0[240][4]}} & loc_sram_buff_w0[240][3:0]) | ({4{loc_sram_buff_w1[240][4]}} & loc_sram_buff_w1[240][3:0]) | ({4{loc_sram_buff_w2[240][4]}} & loc_sram_buff_w2[240][3:0]) | ({4{loc_sram_buff_w3[240][4]}} & loc_sram_buff_w3[240][3:0]) | ({4{loc_sram_buff_w4[240][4]}} & loc_sram_buff_w4[240][3:0]) | ({4{loc_sram_buff_w5[240][4]}} & loc_sram_buff_w5[240][3:0]) | ({4{loc_sram_buff_w6[240][4]}} & loc_sram_buff_w6[240][3:0]) | ({4{loc_sram_buff_w7[240][4]}} & loc_sram_buff_w7[240][3:0]) | ({4{loc_sram_buff_w8[240][4]}} & loc_sram_buff_w8[240][3:0]) | ({4{loc_sram_buff_w9[240][4]}} & loc_sram_buff_w9[240][3:0]) | ({4{loc_sram_buff_w10[240][4]}} & loc_sram_buff_w10[240][3:0]) | ({4{loc_sram_buff_w11[240][4]}} & loc_sram_buff_w11[240][3:0]) | ({4{loc_sram_buff_w12[240][4]}} & loc_sram_buff_w12[240][3:0]) | ({4{loc_sram_buff_w13[240][4]}} & loc_sram_buff_w13[240][3:0]) | ({4{loc_sram_buff_w14[240][4]}} & loc_sram_buff_w14[240][3:0]) | ({4{loc_sram_buff_w15[240][4]}} & loc_sram_buff_w15[240][3:0]);
	loc_rdata_buff[  59:  56] = ({4{loc_sram_buff_w0[241][4]}} & loc_sram_buff_w0[241][3:0]) | ({4{loc_sram_buff_w1[241][4]}} & loc_sram_buff_w1[241][3:0]) | ({4{loc_sram_buff_w2[241][4]}} & loc_sram_buff_w2[241][3:0]) | ({4{loc_sram_buff_w3[241][4]}} & loc_sram_buff_w3[241][3:0]) | ({4{loc_sram_buff_w4[241][4]}} & loc_sram_buff_w4[241][3:0]) | ({4{loc_sram_buff_w5[241][4]}} & loc_sram_buff_w5[241][3:0]) | ({4{loc_sram_buff_w6[241][4]}} & loc_sram_buff_w6[241][3:0]) | ({4{loc_sram_buff_w7[241][4]}} & loc_sram_buff_w7[241][3:0]) | ({4{loc_sram_buff_w8[241][4]}} & loc_sram_buff_w8[241][3:0]) | ({4{loc_sram_buff_w9[241][4]}} & loc_sram_buff_w9[241][3:0]) | ({4{loc_sram_buff_w10[241][4]}} & loc_sram_buff_w10[241][3:0]) | ({4{loc_sram_buff_w11[241][4]}} & loc_sram_buff_w11[241][3:0]) | ({4{loc_sram_buff_w12[241][4]}} & loc_sram_buff_w12[241][3:0]) | ({4{loc_sram_buff_w13[241][4]}} & loc_sram_buff_w13[241][3:0]) | ({4{loc_sram_buff_w14[241][4]}} & loc_sram_buff_w14[241][3:0]) | ({4{loc_sram_buff_w15[241][4]}} & loc_sram_buff_w15[241][3:0]);
	loc_rdata_buff[  55:  52] = ({4{loc_sram_buff_w0[242][4]}} & loc_sram_buff_w0[242][3:0]) | ({4{loc_sram_buff_w1[242][4]}} & loc_sram_buff_w1[242][3:0]) | ({4{loc_sram_buff_w2[242][4]}} & loc_sram_buff_w2[242][3:0]) | ({4{loc_sram_buff_w3[242][4]}} & loc_sram_buff_w3[242][3:0]) | ({4{loc_sram_buff_w4[242][4]}} & loc_sram_buff_w4[242][3:0]) | ({4{loc_sram_buff_w5[242][4]}} & loc_sram_buff_w5[242][3:0]) | ({4{loc_sram_buff_w6[242][4]}} & loc_sram_buff_w6[242][3:0]) | ({4{loc_sram_buff_w7[242][4]}} & loc_sram_buff_w7[242][3:0]) | ({4{loc_sram_buff_w8[242][4]}} & loc_sram_buff_w8[242][3:0]) | ({4{loc_sram_buff_w9[242][4]}} & loc_sram_buff_w9[242][3:0]) | ({4{loc_sram_buff_w10[242][4]}} & loc_sram_buff_w10[242][3:0]) | ({4{loc_sram_buff_w11[242][4]}} & loc_sram_buff_w11[242][3:0]) | ({4{loc_sram_buff_w12[242][4]}} & loc_sram_buff_w12[242][3:0]) | ({4{loc_sram_buff_w13[242][4]}} & loc_sram_buff_w13[242][3:0]) | ({4{loc_sram_buff_w14[242][4]}} & loc_sram_buff_w14[242][3:0]) | ({4{loc_sram_buff_w15[242][4]}} & loc_sram_buff_w15[242][3:0]);
	loc_rdata_buff[  51:  48] = ({4{loc_sram_buff_w0[243][4]}} & loc_sram_buff_w0[243][3:0]) | ({4{loc_sram_buff_w1[243][4]}} & loc_sram_buff_w1[243][3:0]) | ({4{loc_sram_buff_w2[243][4]}} & loc_sram_buff_w2[243][3:0]) | ({4{loc_sram_buff_w3[243][4]}} & loc_sram_buff_w3[243][3:0]) | ({4{loc_sram_buff_w4[243][4]}} & loc_sram_buff_w4[243][3:0]) | ({4{loc_sram_buff_w5[243][4]}} & loc_sram_buff_w5[243][3:0]) | ({4{loc_sram_buff_w6[243][4]}} & loc_sram_buff_w6[243][3:0]) | ({4{loc_sram_buff_w7[243][4]}} & loc_sram_buff_w7[243][3:0]) | ({4{loc_sram_buff_w8[243][4]}} & loc_sram_buff_w8[243][3:0]) | ({4{loc_sram_buff_w9[243][4]}} & loc_sram_buff_w9[243][3:0]) | ({4{loc_sram_buff_w10[243][4]}} & loc_sram_buff_w10[243][3:0]) | ({4{loc_sram_buff_w11[243][4]}} & loc_sram_buff_w11[243][3:0]) | ({4{loc_sram_buff_w12[243][4]}} & loc_sram_buff_w12[243][3:0]) | ({4{loc_sram_buff_w13[243][4]}} & loc_sram_buff_w13[243][3:0]) | ({4{loc_sram_buff_w14[243][4]}} & loc_sram_buff_w14[243][3:0]) | ({4{loc_sram_buff_w15[243][4]}} & loc_sram_buff_w15[243][3:0]);
	loc_rdata_buff[  47:  44] = ({4{loc_sram_buff_w0[244][4]}} & loc_sram_buff_w0[244][3:0]) | ({4{loc_sram_buff_w1[244][4]}} & loc_sram_buff_w1[244][3:0]) | ({4{loc_sram_buff_w2[244][4]}} & loc_sram_buff_w2[244][3:0]) | ({4{loc_sram_buff_w3[244][4]}} & loc_sram_buff_w3[244][3:0]) | ({4{loc_sram_buff_w4[244][4]}} & loc_sram_buff_w4[244][3:0]) | ({4{loc_sram_buff_w5[244][4]}} & loc_sram_buff_w5[244][3:0]) | ({4{loc_sram_buff_w6[244][4]}} & loc_sram_buff_w6[244][3:0]) | ({4{loc_sram_buff_w7[244][4]}} & loc_sram_buff_w7[244][3:0]) | ({4{loc_sram_buff_w8[244][4]}} & loc_sram_buff_w8[244][3:0]) | ({4{loc_sram_buff_w9[244][4]}} & loc_sram_buff_w9[244][3:0]) | ({4{loc_sram_buff_w10[244][4]}} & loc_sram_buff_w10[244][3:0]) | ({4{loc_sram_buff_w11[244][4]}} & loc_sram_buff_w11[244][3:0]) | ({4{loc_sram_buff_w12[244][4]}} & loc_sram_buff_w12[244][3:0]) | ({4{loc_sram_buff_w13[244][4]}} & loc_sram_buff_w13[244][3:0]) | ({4{loc_sram_buff_w14[244][4]}} & loc_sram_buff_w14[244][3:0]) | ({4{loc_sram_buff_w15[244][4]}} & loc_sram_buff_w15[244][3:0]);
	loc_rdata_buff[  43:  40] = ({4{loc_sram_buff_w0[245][4]}} & loc_sram_buff_w0[245][3:0]) | ({4{loc_sram_buff_w1[245][4]}} & loc_sram_buff_w1[245][3:0]) | ({4{loc_sram_buff_w2[245][4]}} & loc_sram_buff_w2[245][3:0]) | ({4{loc_sram_buff_w3[245][4]}} & loc_sram_buff_w3[245][3:0]) | ({4{loc_sram_buff_w4[245][4]}} & loc_sram_buff_w4[245][3:0]) | ({4{loc_sram_buff_w5[245][4]}} & loc_sram_buff_w5[245][3:0]) | ({4{loc_sram_buff_w6[245][4]}} & loc_sram_buff_w6[245][3:0]) | ({4{loc_sram_buff_w7[245][4]}} & loc_sram_buff_w7[245][3:0]) | ({4{loc_sram_buff_w8[245][4]}} & loc_sram_buff_w8[245][3:0]) | ({4{loc_sram_buff_w9[245][4]}} & loc_sram_buff_w9[245][3:0]) | ({4{loc_sram_buff_w10[245][4]}} & loc_sram_buff_w10[245][3:0]) | ({4{loc_sram_buff_w11[245][4]}} & loc_sram_buff_w11[245][3:0]) | ({4{loc_sram_buff_w12[245][4]}} & loc_sram_buff_w12[245][3:0]) | ({4{loc_sram_buff_w13[245][4]}} & loc_sram_buff_w13[245][3:0]) | ({4{loc_sram_buff_w14[245][4]}} & loc_sram_buff_w14[245][3:0]) | ({4{loc_sram_buff_w15[245][4]}} & loc_sram_buff_w15[245][3:0]);
	loc_rdata_buff[  39:  36] = ({4{loc_sram_buff_w0[246][4]}} & loc_sram_buff_w0[246][3:0]) | ({4{loc_sram_buff_w1[246][4]}} & loc_sram_buff_w1[246][3:0]) | ({4{loc_sram_buff_w2[246][4]}} & loc_sram_buff_w2[246][3:0]) | ({4{loc_sram_buff_w3[246][4]}} & loc_sram_buff_w3[246][3:0]) | ({4{loc_sram_buff_w4[246][4]}} & loc_sram_buff_w4[246][3:0]) | ({4{loc_sram_buff_w5[246][4]}} & loc_sram_buff_w5[246][3:0]) | ({4{loc_sram_buff_w6[246][4]}} & loc_sram_buff_w6[246][3:0]) | ({4{loc_sram_buff_w7[246][4]}} & loc_sram_buff_w7[246][3:0]) | ({4{loc_sram_buff_w8[246][4]}} & loc_sram_buff_w8[246][3:0]) | ({4{loc_sram_buff_w9[246][4]}} & loc_sram_buff_w9[246][3:0]) | ({4{loc_sram_buff_w10[246][4]}} & loc_sram_buff_w10[246][3:0]) | ({4{loc_sram_buff_w11[246][4]}} & loc_sram_buff_w11[246][3:0]) | ({4{loc_sram_buff_w12[246][4]}} & loc_sram_buff_w12[246][3:0]) | ({4{loc_sram_buff_w13[246][4]}} & loc_sram_buff_w13[246][3:0]) | ({4{loc_sram_buff_w14[246][4]}} & loc_sram_buff_w14[246][3:0]) | ({4{loc_sram_buff_w15[246][4]}} & loc_sram_buff_w15[246][3:0]);
	loc_rdata_buff[  35:  32] = ({4{loc_sram_buff_w0[247][4]}} & loc_sram_buff_w0[247][3:0]) | ({4{loc_sram_buff_w1[247][4]}} & loc_sram_buff_w1[247][3:0]) | ({4{loc_sram_buff_w2[247][4]}} & loc_sram_buff_w2[247][3:0]) | ({4{loc_sram_buff_w3[247][4]}} & loc_sram_buff_w3[247][3:0]) | ({4{loc_sram_buff_w4[247][4]}} & loc_sram_buff_w4[247][3:0]) | ({4{loc_sram_buff_w5[247][4]}} & loc_sram_buff_w5[247][3:0]) | ({4{loc_sram_buff_w6[247][4]}} & loc_sram_buff_w6[247][3:0]) | ({4{loc_sram_buff_w7[247][4]}} & loc_sram_buff_w7[247][3:0]) | ({4{loc_sram_buff_w8[247][4]}} & loc_sram_buff_w8[247][3:0]) | ({4{loc_sram_buff_w9[247][4]}} & loc_sram_buff_w9[247][3:0]) | ({4{loc_sram_buff_w10[247][4]}} & loc_sram_buff_w10[247][3:0]) | ({4{loc_sram_buff_w11[247][4]}} & loc_sram_buff_w11[247][3:0]) | ({4{loc_sram_buff_w12[247][4]}} & loc_sram_buff_w12[247][3:0]) | ({4{loc_sram_buff_w13[247][4]}} & loc_sram_buff_w13[247][3:0]) | ({4{loc_sram_buff_w14[247][4]}} & loc_sram_buff_w14[247][3:0]) | ({4{loc_sram_buff_w15[247][4]}} & loc_sram_buff_w15[247][3:0]);
	loc_rdata_buff[  31:  28] = ({4{loc_sram_buff_w0[248][4]}} & loc_sram_buff_w0[248][3:0]) | ({4{loc_sram_buff_w1[248][4]}} & loc_sram_buff_w1[248][3:0]) | ({4{loc_sram_buff_w2[248][4]}} & loc_sram_buff_w2[248][3:0]) | ({4{loc_sram_buff_w3[248][4]}} & loc_sram_buff_w3[248][3:0]) | ({4{loc_sram_buff_w4[248][4]}} & loc_sram_buff_w4[248][3:0]) | ({4{loc_sram_buff_w5[248][4]}} & loc_sram_buff_w5[248][3:0]) | ({4{loc_sram_buff_w6[248][4]}} & loc_sram_buff_w6[248][3:0]) | ({4{loc_sram_buff_w7[248][4]}} & loc_sram_buff_w7[248][3:0]) | ({4{loc_sram_buff_w8[248][4]}} & loc_sram_buff_w8[248][3:0]) | ({4{loc_sram_buff_w9[248][4]}} & loc_sram_buff_w9[248][3:0]) | ({4{loc_sram_buff_w10[248][4]}} & loc_sram_buff_w10[248][3:0]) | ({4{loc_sram_buff_w11[248][4]}} & loc_sram_buff_w11[248][3:0]) | ({4{loc_sram_buff_w12[248][4]}} & loc_sram_buff_w12[248][3:0]) | ({4{loc_sram_buff_w13[248][4]}} & loc_sram_buff_w13[248][3:0]) | ({4{loc_sram_buff_w14[248][4]}} & loc_sram_buff_w14[248][3:0]) | ({4{loc_sram_buff_w15[248][4]}} & loc_sram_buff_w15[248][3:0]);
	loc_rdata_buff[  27:  24] = ({4{loc_sram_buff_w0[249][4]}} & loc_sram_buff_w0[249][3:0]) | ({4{loc_sram_buff_w1[249][4]}} & loc_sram_buff_w1[249][3:0]) | ({4{loc_sram_buff_w2[249][4]}} & loc_sram_buff_w2[249][3:0]) | ({4{loc_sram_buff_w3[249][4]}} & loc_sram_buff_w3[249][3:0]) | ({4{loc_sram_buff_w4[249][4]}} & loc_sram_buff_w4[249][3:0]) | ({4{loc_sram_buff_w5[249][4]}} & loc_sram_buff_w5[249][3:0]) | ({4{loc_sram_buff_w6[249][4]}} & loc_sram_buff_w6[249][3:0]) | ({4{loc_sram_buff_w7[249][4]}} & loc_sram_buff_w7[249][3:0]) | ({4{loc_sram_buff_w8[249][4]}} & loc_sram_buff_w8[249][3:0]) | ({4{loc_sram_buff_w9[249][4]}} & loc_sram_buff_w9[249][3:0]) | ({4{loc_sram_buff_w10[249][4]}} & loc_sram_buff_w10[249][3:0]) | ({4{loc_sram_buff_w11[249][4]}} & loc_sram_buff_w11[249][3:0]) | ({4{loc_sram_buff_w12[249][4]}} & loc_sram_buff_w12[249][3:0]) | ({4{loc_sram_buff_w13[249][4]}} & loc_sram_buff_w13[249][3:0]) | ({4{loc_sram_buff_w14[249][4]}} & loc_sram_buff_w14[249][3:0]) | ({4{loc_sram_buff_w15[249][4]}} & loc_sram_buff_w15[249][3:0]);
	loc_rdata_buff[  23:  20] = ({4{loc_sram_buff_w0[250][4]}} & loc_sram_buff_w0[250][3:0]) | ({4{loc_sram_buff_w1[250][4]}} & loc_sram_buff_w1[250][3:0]) | ({4{loc_sram_buff_w2[250][4]}} & loc_sram_buff_w2[250][3:0]) | ({4{loc_sram_buff_w3[250][4]}} & loc_sram_buff_w3[250][3:0]) | ({4{loc_sram_buff_w4[250][4]}} & loc_sram_buff_w4[250][3:0]) | ({4{loc_sram_buff_w5[250][4]}} & loc_sram_buff_w5[250][3:0]) | ({4{loc_sram_buff_w6[250][4]}} & loc_sram_buff_w6[250][3:0]) | ({4{loc_sram_buff_w7[250][4]}} & loc_sram_buff_w7[250][3:0]) | ({4{loc_sram_buff_w8[250][4]}} & loc_sram_buff_w8[250][3:0]) | ({4{loc_sram_buff_w9[250][4]}} & loc_sram_buff_w9[250][3:0]) | ({4{loc_sram_buff_w10[250][4]}} & loc_sram_buff_w10[250][3:0]) | ({4{loc_sram_buff_w11[250][4]}} & loc_sram_buff_w11[250][3:0]) | ({4{loc_sram_buff_w12[250][4]}} & loc_sram_buff_w12[250][3:0]) | ({4{loc_sram_buff_w13[250][4]}} & loc_sram_buff_w13[250][3:0]) | ({4{loc_sram_buff_w14[250][4]}} & loc_sram_buff_w14[250][3:0]) | ({4{loc_sram_buff_w15[250][4]}} & loc_sram_buff_w15[250][3:0]);
	loc_rdata_buff[  19:  16] = ({4{loc_sram_buff_w0[251][4]}} & loc_sram_buff_w0[251][3:0]) | ({4{loc_sram_buff_w1[251][4]}} & loc_sram_buff_w1[251][3:0]) | ({4{loc_sram_buff_w2[251][4]}} & loc_sram_buff_w2[251][3:0]) | ({4{loc_sram_buff_w3[251][4]}} & loc_sram_buff_w3[251][3:0]) | ({4{loc_sram_buff_w4[251][4]}} & loc_sram_buff_w4[251][3:0]) | ({4{loc_sram_buff_w5[251][4]}} & loc_sram_buff_w5[251][3:0]) | ({4{loc_sram_buff_w6[251][4]}} & loc_sram_buff_w6[251][3:0]) | ({4{loc_sram_buff_w7[251][4]}} & loc_sram_buff_w7[251][3:0]) | ({4{loc_sram_buff_w8[251][4]}} & loc_sram_buff_w8[251][3:0]) | ({4{loc_sram_buff_w9[251][4]}} & loc_sram_buff_w9[251][3:0]) | ({4{loc_sram_buff_w10[251][4]}} & loc_sram_buff_w10[251][3:0]) | ({4{loc_sram_buff_w11[251][4]}} & loc_sram_buff_w11[251][3:0]) | ({4{loc_sram_buff_w12[251][4]}} & loc_sram_buff_w12[251][3:0]) | ({4{loc_sram_buff_w13[251][4]}} & loc_sram_buff_w13[251][3:0]) | ({4{loc_sram_buff_w14[251][4]}} & loc_sram_buff_w14[251][3:0]) | ({4{loc_sram_buff_w15[251][4]}} & loc_sram_buff_w15[251][3:0]);
	loc_rdata_buff[  15:  12] = ({4{loc_sram_buff_w0[252][4]}} & loc_sram_buff_w0[252][3:0]) | ({4{loc_sram_buff_w1[252][4]}} & loc_sram_buff_w1[252][3:0]) | ({4{loc_sram_buff_w2[252][4]}} & loc_sram_buff_w2[252][3:0]) | ({4{loc_sram_buff_w3[252][4]}} & loc_sram_buff_w3[252][3:0]) | ({4{loc_sram_buff_w4[252][4]}} & loc_sram_buff_w4[252][3:0]) | ({4{loc_sram_buff_w5[252][4]}} & loc_sram_buff_w5[252][3:0]) | ({4{loc_sram_buff_w6[252][4]}} & loc_sram_buff_w6[252][3:0]) | ({4{loc_sram_buff_w7[252][4]}} & loc_sram_buff_w7[252][3:0]) | ({4{loc_sram_buff_w8[252][4]}} & loc_sram_buff_w8[252][3:0]) | ({4{loc_sram_buff_w9[252][4]}} & loc_sram_buff_w9[252][3:0]) | ({4{loc_sram_buff_w10[252][4]}} & loc_sram_buff_w10[252][3:0]) | ({4{loc_sram_buff_w11[252][4]}} & loc_sram_buff_w11[252][3:0]) | ({4{loc_sram_buff_w12[252][4]}} & loc_sram_buff_w12[252][3:0]) | ({4{loc_sram_buff_w13[252][4]}} & loc_sram_buff_w13[252][3:0]) | ({4{loc_sram_buff_w14[252][4]}} & loc_sram_buff_w14[252][3:0]) | ({4{loc_sram_buff_w15[252][4]}} & loc_sram_buff_w15[252][3:0]);
	loc_rdata_buff[  11:   8] = ({4{loc_sram_buff_w0[253][4]}} & loc_sram_buff_w0[253][3:0]) | ({4{loc_sram_buff_w1[253][4]}} & loc_sram_buff_w1[253][3:0]) | ({4{loc_sram_buff_w2[253][4]}} & loc_sram_buff_w2[253][3:0]) | ({4{loc_sram_buff_w3[253][4]}} & loc_sram_buff_w3[253][3:0]) | ({4{loc_sram_buff_w4[253][4]}} & loc_sram_buff_w4[253][3:0]) | ({4{loc_sram_buff_w5[253][4]}} & loc_sram_buff_w5[253][3:0]) | ({4{loc_sram_buff_w6[253][4]}} & loc_sram_buff_w6[253][3:0]) | ({4{loc_sram_buff_w7[253][4]}} & loc_sram_buff_w7[253][3:0]) | ({4{loc_sram_buff_w8[253][4]}} & loc_sram_buff_w8[253][3:0]) | ({4{loc_sram_buff_w9[253][4]}} & loc_sram_buff_w9[253][3:0]) | ({4{loc_sram_buff_w10[253][4]}} & loc_sram_buff_w10[253][3:0]) | ({4{loc_sram_buff_w11[253][4]}} & loc_sram_buff_w11[253][3:0]) | ({4{loc_sram_buff_w12[253][4]}} & loc_sram_buff_w12[253][3:0]) | ({4{loc_sram_buff_w13[253][4]}} & loc_sram_buff_w13[253][3:0]) | ({4{loc_sram_buff_w14[253][4]}} & loc_sram_buff_w14[253][3:0]) | ({4{loc_sram_buff_w15[253][4]}} & loc_sram_buff_w15[253][3:0]);
	loc_rdata_buff[   7:   4] = ({4{loc_sram_buff_w0[254][4]}} & loc_sram_buff_w0[254][3:0]) | ({4{loc_sram_buff_w1[254][4]}} & loc_sram_buff_w1[254][3:0]) | ({4{loc_sram_buff_w2[254][4]}} & loc_sram_buff_w2[254][3:0]) | ({4{loc_sram_buff_w3[254][4]}} & loc_sram_buff_w3[254][3:0]) | ({4{loc_sram_buff_w4[254][4]}} & loc_sram_buff_w4[254][3:0]) | ({4{loc_sram_buff_w5[254][4]}} & loc_sram_buff_w5[254][3:0]) | ({4{loc_sram_buff_w6[254][4]}} & loc_sram_buff_w6[254][3:0]) | ({4{loc_sram_buff_w7[254][4]}} & loc_sram_buff_w7[254][3:0]) | ({4{loc_sram_buff_w8[254][4]}} & loc_sram_buff_w8[254][3:0]) | ({4{loc_sram_buff_w9[254][4]}} & loc_sram_buff_w9[254][3:0]) | ({4{loc_sram_buff_w10[254][4]}} & loc_sram_buff_w10[254][3:0]) | ({4{loc_sram_buff_w11[254][4]}} & loc_sram_buff_w11[254][3:0]) | ({4{loc_sram_buff_w12[254][4]}} & loc_sram_buff_w12[254][3:0]) | ({4{loc_sram_buff_w13[254][4]}} & loc_sram_buff_w13[254][3:0]) | ({4{loc_sram_buff_w14[254][4]}} & loc_sram_buff_w14[254][3:0]) | ({4{loc_sram_buff_w15[254][4]}} & loc_sram_buff_w15[254][3:0]);
	loc_rdata_buff[   3:   0] = ({4{loc_sram_buff_w0[255][4]}} & loc_sram_buff_w0[255][3:0]) | ({4{loc_sram_buff_w1[255][4]}} & loc_sram_buff_w1[255][3:0]) | ({4{loc_sram_buff_w2[255][4]}} & loc_sram_buff_w2[255][3:0]) | ({4{loc_sram_buff_w3[255][4]}} & loc_sram_buff_w3[255][3:0]) | ({4{loc_sram_buff_w4[255][4]}} & loc_sram_buff_w4[255][3:0]) | ({4{loc_sram_buff_w5[255][4]}} & loc_sram_buff_w5[255][3:0]) | ({4{loc_sram_buff_w6[255][4]}} & loc_sram_buff_w6[255][3:0]) | ({4{loc_sram_buff_w7[255][4]}} & loc_sram_buff_w7[255][3:0]) | ({4{loc_sram_buff_w8[255][4]}} & loc_sram_buff_w8[255][3:0]) | ({4{loc_sram_buff_w9[255][4]}} & loc_sram_buff_w9[255][3:0]) | ({4{loc_sram_buff_w10[255][4]}} & loc_sram_buff_w10[255][3:0]) | ({4{loc_sram_buff_w11[255][4]}} & loc_sram_buff_w11[255][3:0]) | ({4{loc_sram_buff_w12[255][4]}} & loc_sram_buff_w12[255][3:0]) | ({4{loc_sram_buff_w13[255][4]}} & loc_sram_buff_w13[255][3:0]) | ({4{loc_sram_buff_w14[255][4]}} & loc_sram_buff_w14[255][3:0]) | ({4{loc_sram_buff_w15[255][4]}} & loc_sram_buff_w15[255][3:0]);

end 

assign w0_loc_rdata = loc_rdata_buff;
assign w1_loc_rdata = loc_rdata_buff;
assign w2_loc_rdata = loc_rdata_buff;
assign w3_loc_rdata = loc_rdata_buff;
assign w4_loc_rdata = loc_rdata_buff;
assign w5_loc_rdata = loc_rdata_buff;
assign w6_loc_rdata = loc_rdata_buff;
assign w7_loc_rdata = loc_rdata_buff;
assign w8_loc_rdata = loc_rdata_buff;
assign w9_loc_rdata = loc_rdata_buff;
assign w10_loc_rdata = loc_rdata_buff;
assign w11_loc_rdata = loc_rdata_buff;
assign w12_loc_rdata = loc_rdata_buff;
assign w13_loc_rdata = loc_rdata_buff;
assign w14_loc_rdata = loc_rdata_buff;
assign w15_loc_rdata = loc_rdata_buff;


always @* begin
	(* synthesis, parallel_case *)
	case(epoch_buff[7:4])
		4'd0: in_mi_j  = {w0_proposal_num0,w0_proposal_num1,w0_proposal_num2,w0_proposal_num3,w0_proposal_num4,w0_proposal_num5,w0_proposal_num6,w0_proposal_num7,w0_proposal_num8,w0_proposal_num9,w0_proposal_num10,w0_proposal_num11,w0_proposal_num12,w0_proposal_num13,w0_proposal_num14,w0_proposal_num15};
	    4'd1: in_mi_j  = {w1_proposal_num0,w1_proposal_num1,w1_proposal_num2,w1_proposal_num3,w1_proposal_num4,w1_proposal_num5,w1_proposal_num6,w1_proposal_num7,w1_proposal_num8,w1_proposal_num9,w1_proposal_num10,w1_proposal_num11,w1_proposal_num12,w1_proposal_num13,w1_proposal_num14,w1_proposal_num15};
	    4'd2: in_mi_j  = {w2_proposal_num0,w2_proposal_num1,w2_proposal_num2,w2_proposal_num3,w2_proposal_num4,w2_proposal_num5,w2_proposal_num6,w2_proposal_num7,w2_proposal_num8,w2_proposal_num9,w2_proposal_num10,w2_proposal_num11,w2_proposal_num12,w2_proposal_num13,w2_proposal_num14,w2_proposal_num15};
	    4'd3: in_mi_j  = {w3_proposal_num0,w3_proposal_num1,w3_proposal_num2,w3_proposal_num3,w3_proposal_num4,w3_proposal_num5,w3_proposal_num6,w3_proposal_num7,w3_proposal_num8,w3_proposal_num9,w3_proposal_num10,w3_proposal_num11,w3_proposal_num12,w3_proposal_num13,w3_proposal_num14,w3_proposal_num15};
	    4'd4: in_mi_j  = {w4_proposal_num0,w4_proposal_num1,w4_proposal_num2,w4_proposal_num3,w4_proposal_num4,w4_proposal_num5,w4_proposal_num6,w4_proposal_num7,w4_proposal_num8,w4_proposal_num9,w4_proposal_num10,w4_proposal_num11,w4_proposal_num12,w4_proposal_num13,w4_proposal_num14,w4_proposal_num15};
	    4'd5: in_mi_j  = {w5_proposal_num0,w5_proposal_num1,w5_proposal_num2,w5_proposal_num3,w5_proposal_num4,w5_proposal_num5,w5_proposal_num6,w5_proposal_num7,w5_proposal_num8,w5_proposal_num9,w5_proposal_num10,w5_proposal_num11,w5_proposal_num12,w5_proposal_num13,w5_proposal_num14,w5_proposal_num15};
	   	4'd6: in_mi_j  = {w6_proposal_num0,w6_proposal_num1,w6_proposal_num2,w6_proposal_num3,w6_proposal_num4,w6_proposal_num5,w6_proposal_num6,w6_proposal_num7,w6_proposal_num8,w6_proposal_num9,w6_proposal_num10,w6_proposal_num11,w6_proposal_num12,w6_proposal_num13,w6_proposal_num14,w6_proposal_num15};
	   	4'd7: in_mi_j  = {w7_proposal_num0,w7_proposal_num1,w7_proposal_num2,w7_proposal_num3,w7_proposal_num4,w7_proposal_num5,w7_proposal_num6,w7_proposal_num7,w7_proposal_num8,w7_proposal_num9,w7_proposal_num10,w7_proposal_num11,w7_proposal_num12,w7_proposal_num13,w7_proposal_num14,w7_proposal_num15};
	   	4'd8: in_mi_j  = {w8_proposal_num0,w8_proposal_num1,w8_proposal_num2,w8_proposal_num3,w8_proposal_num4,w8_proposal_num5,w8_proposal_num6,w8_proposal_num7,w8_proposal_num8,w8_proposal_num9,w8_proposal_num10,w8_proposal_num11,w8_proposal_num12,w8_proposal_num13,w8_proposal_num14,w8_proposal_num15};
	   	4'd9: in_mi_j  = {w9_proposal_num0,w9_proposal_num1,w9_proposal_num2,w9_proposal_num3,w9_proposal_num4,w9_proposal_num5,w9_proposal_num6,w9_proposal_num7,w9_proposal_num8,w9_proposal_num9,w9_proposal_num10,w9_proposal_num11,w9_proposal_num12,w9_proposal_num13,w9_proposal_num14,w9_proposal_num15};
	   	4'd10: in_mi_j = {w10_proposal_num0,w10_proposal_num1,w10_proposal_num2,w10_proposal_num3,w10_proposal_num4,w10_proposal_num5,w10_proposal_num6,w10_proposal_num7,w10_proposal_num8,w10_proposal_num9,w10_proposal_num10,w10_proposal_num11,w10_proposal_num12,w10_proposal_num13,w10_proposal_num14,w10_proposal_num15};
	   	4'd11: in_mi_j = {w11_proposal_num0,w11_proposal_num1,w11_proposal_num2,w11_proposal_num3,w11_proposal_num4,w11_proposal_num5,w11_proposal_num6,w11_proposal_num7,w11_proposal_num8,w11_proposal_num9,w11_proposal_num10,w11_proposal_num11,w11_proposal_num12,w11_proposal_num13,w11_proposal_num14,w11_proposal_num15};
		4'd12: in_mi_j = {w12_proposal_num0,w12_proposal_num1,w12_proposal_num2,w12_proposal_num3,w12_proposal_num4,w12_proposal_num5,w12_proposal_num6,w12_proposal_num7,w12_proposal_num8,w12_proposal_num9,w12_proposal_num10,w12_proposal_num11,w12_proposal_num12,w12_proposal_num13,w12_proposal_num14,w12_proposal_num15};
	   	4'd13: in_mi_j = {w13_proposal_num0,w13_proposal_num1,w13_proposal_num2,w13_proposal_num3,w13_proposal_num4,w13_proposal_num5,w13_proposal_num6,w13_proposal_num7,w13_proposal_num8,w13_proposal_num9,w13_proposal_num10,w13_proposal_num11,w13_proposal_num12,w13_proposal_num13,w13_proposal_num14,w13_proposal_num15};
	   	4'd14: in_mi_j = {w14_proposal_num0,w14_proposal_num1,w14_proposal_num2,w14_proposal_num3,w14_proposal_num4,w14_proposal_num5,w14_proposal_num6,w14_proposal_num7,w14_proposal_num8,w14_proposal_num9,w14_proposal_num10,w14_proposal_num11,w14_proposal_num12,w14_proposal_num13,w14_proposal_num14,w14_proposal_num15};
	   	4'd15: in_mi_j = {w15_proposal_num0,w15_proposal_num1,w15_proposal_num2,w15_proposal_num3,w15_proposal_num4,w15_proposal_num5,w15_proposal_num6,w15_proposal_num7,w15_proposal_num8,w15_proposal_num9,w15_proposal_num10,w15_proposal_num11,w15_proposal_num12,w15_proposal_num13,w15_proposal_num14,w15_proposal_num15};
	endcase 

	(* synthesis, parallel_case *)
	case(epoch_buff[7:4]) 
	4'd0:	in_mj_i = {w0_proposal_num0,w1_proposal_num0,w2_proposal_num0,w3_proposal_num0,w4_proposal_num0,w5_proposal_num0,w6_proposal_num0,w7_proposal_num0,w8_proposal_num0,w9_proposal_num0,w10_proposal_num0,w11_proposal_num0,w12_proposal_num0,w13_proposal_num0,w14_proposal_num0,w15_proposal_num0};
	4'd1:	in_mj_i = {w0_proposal_num1,w1_proposal_num1,w2_proposal_num1,w3_proposal_num1,w4_proposal_num1,w5_proposal_num1,w6_proposal_num1,w7_proposal_num1,w8_proposal_num1,w9_proposal_num1,w10_proposal_num1,w11_proposal_num1,w12_proposal_num1,w13_proposal_num1,w14_proposal_num1,w15_proposal_num1};
	4'd2:	in_mj_i = {w0_proposal_num2,w1_proposal_num2,w2_proposal_num2,w3_proposal_num2,w4_proposal_num2,w5_proposal_num2,w6_proposal_num2,w7_proposal_num2,w8_proposal_num2,w9_proposal_num2,w10_proposal_num2,w11_proposal_num2,w12_proposal_num2,w13_proposal_num2,w14_proposal_num2,w15_proposal_num2};
	4'd3:	in_mj_i = {w0_proposal_num3,w1_proposal_num3,w2_proposal_num3,w3_proposal_num3,w4_proposal_num3,w5_proposal_num3,w6_proposal_num3,w7_proposal_num3,w8_proposal_num3,w9_proposal_num3,w10_proposal_num3,w11_proposal_num3,w12_proposal_num3,w13_proposal_num3,w14_proposal_num3,w15_proposal_num3};
	4'd4:	in_mj_i = {w0_proposal_num4,w1_proposal_num4,w2_proposal_num4,w3_proposal_num4,w4_proposal_num4,w5_proposal_num4,w6_proposal_num4,w7_proposal_num4,w8_proposal_num4,w9_proposal_num4,w10_proposal_num4,w11_proposal_num4,w12_proposal_num4,w13_proposal_num4,w14_proposal_num4,w15_proposal_num4};
	4'd5:	in_mj_i = {w0_proposal_num5,w1_proposal_num5,w2_proposal_num5,w3_proposal_num5,w4_proposal_num5,w5_proposal_num5,w6_proposal_num5,w7_proposal_num5,w8_proposal_num5,w9_proposal_num5,w10_proposal_num5,w11_proposal_num5,w12_proposal_num5,w13_proposal_num5,w14_proposal_num5,w15_proposal_num5};
	4'd6:	in_mj_i = {w0_proposal_num6,w1_proposal_num6,w2_proposal_num6,w3_proposal_num6,w4_proposal_num6,w5_proposal_num6,w6_proposal_num6,w7_proposal_num6,w8_proposal_num6,w9_proposal_num6,w10_proposal_num6,w11_proposal_num6,w12_proposal_num6,w13_proposal_num6,w14_proposal_num6,w15_proposal_num6};
	4'd7:	in_mj_i = {w0_proposal_num7,w1_proposal_num7,w2_proposal_num7,w3_proposal_num7,w4_proposal_num7,w5_proposal_num7,w6_proposal_num7,w7_proposal_num7,w8_proposal_num7,w9_proposal_num7,w10_proposal_num7,w11_proposal_num7,w12_proposal_num7,w13_proposal_num7,w14_proposal_num7,w15_proposal_num7};
	4'd8:	in_mj_i = {w0_proposal_num8,w1_proposal_num8,w2_proposal_num8,w3_proposal_num8,w4_proposal_num8,w5_proposal_num8,w6_proposal_num8,w7_proposal_num8,w8_proposal_num8,w9_proposal_num8,w10_proposal_num8,w11_proposal_num8,w12_proposal_num8,w13_proposal_num8,w14_proposal_num8,w15_proposal_num8};
	4'd9:	in_mj_i = {w0_proposal_num9,w1_proposal_num9,w2_proposal_num9,w3_proposal_num9,w4_proposal_num9,w5_proposal_num9,w6_proposal_num9,w7_proposal_num9,w8_proposal_num9,w9_proposal_num9,w10_proposal_num9,w11_proposal_num9,w12_proposal_num9,w13_proposal_num9,w14_proposal_num9,w15_proposal_num9};
	4'd10:	in_mj_i = {w0_proposal_num10,w1_proposal_num10,w2_proposal_num10,w3_proposal_num10,w4_proposal_num10,w5_proposal_num10,w6_proposal_num10,w7_proposal_num10,w8_proposal_num10,w9_proposal_num10,w10_proposal_num10,w11_proposal_num10,w12_proposal_num10,w13_proposal_num10,w14_proposal_num10,w15_proposal_num10};
	4'd11:	in_mj_i = {w0_proposal_num11,w1_proposal_num11,w2_proposal_num11,w3_proposal_num11,w4_proposal_num11,w5_proposal_num11,w6_proposal_num11,w7_proposal_num11,w8_proposal_num11,w9_proposal_num11,w10_proposal_num11,w11_proposal_num11,w12_proposal_num11,w13_proposal_num11,w14_proposal_num11,w15_proposal_num11};
	4'd12:	in_mj_i = {w0_proposal_num12,w1_proposal_num12,w2_proposal_num12,w3_proposal_num12,w4_proposal_num12,w5_proposal_num12,w6_proposal_num12,w7_proposal_num12,w8_proposal_num12,w9_proposal_num12,w10_proposal_num12,w11_proposal_num12,w12_proposal_num12,w13_proposal_num12,w14_proposal_num12,w15_proposal_num12};
	4'd13:	in_mj_i = {w0_proposal_num13,w1_proposal_num13,w2_proposal_num13,w3_proposal_num13,w4_proposal_num13,w5_proposal_num13,w6_proposal_num13,w7_proposal_num13,w8_proposal_num13,w9_proposal_num13,w10_proposal_num13,w11_proposal_num13,w12_proposal_num13,w13_proposal_num13,w14_proposal_num13,w15_proposal_num13};
	4'd14:	in_mj_i = {w0_proposal_num14,w1_proposal_num14,w2_proposal_num14,w3_proposal_num14,w4_proposal_num14,w5_proposal_num14,w6_proposal_num14,w7_proposal_num14,w8_proposal_num14,w9_proposal_num14,w10_proposal_num14,w11_proposal_num14,w12_proposal_num14,w13_proposal_num14,w14_proposal_num14,w15_proposal_num14};
	4'd15:	in_mj_i = {w0_proposal_num15,w1_proposal_num15,w2_proposal_num15,w3_proposal_num15,w4_proposal_num15,w5_proposal_num15,w6_proposal_num15,w7_proposal_num15,w8_proposal_num15,w9_proposal_num15,w10_proposal_num15,w11_proposal_num15,w12_proposal_num15,w13_proposal_num15,w14_proposal_num15,w15_proposal_num15};
		
	endcase 
end 

// vid sram read in
always @* begin 
	if(state <= WORKER) begin 
		vid_sram_raddr0 = {iter[0], batch_num[7:4]};	vid_sram_raddr8 = {iter[0], batch_num[7:4]};
		vid_sram_raddr1 = {iter[0], batch_num[7:4]};	vid_sram_raddr9 = {iter[0], batch_num[7:4]};
		vid_sram_raddr2 = {iter[0], batch_num[7:4]};	vid_sram_raddr10 = {iter[0], batch_num[7:4]};
		vid_sram_raddr3 = {iter[0], batch_num[7:4]};	vid_sram_raddr11 = {iter[0], batch_num[7:4]};
		vid_sram_raddr4 = {iter[0], batch_num[7:4]};	vid_sram_raddr12 = {iter[0], batch_num[7:4]};
		vid_sram_raddr5 = {iter[0], batch_num[7:4]};	vid_sram_raddr13 = {iter[0], batch_num[7:4]};
		vid_sram_raddr6 = {iter[0], batch_num[7:4]};	vid_sram_raddr14 = {iter[0], batch_num[7:4]};
		vid_sram_raddr7 = {iter[0], batch_num[7:4]};	vid_sram_raddr15 = {iter[0], batch_num[7:4]};
	end else begin 
		vid_sram_raddr0 = vid_sram_raddr_total; vid_sram_raddr8 = vid_sram_raddr_total;
		vid_sram_raddr1 = vid_sram_raddr_total; vid_sram_raddr9 = vid_sram_raddr_total;
		vid_sram_raddr2 = vid_sram_raddr_total; vid_sram_raddr10 = vid_sram_raddr_total;
		vid_sram_raddr3 = vid_sram_raddr_total; vid_sram_raddr11 = vid_sram_raddr_total;
		vid_sram_raddr4 = vid_sram_raddr_total; vid_sram_raddr12 = vid_sram_raddr_total;
		vid_sram_raddr5 = vid_sram_raddr_total; vid_sram_raddr13 = vid_sram_raddr_total;
		vid_sram_raddr6 = vid_sram_raddr_total; vid_sram_raddr14 = vid_sram_raddr_total;
		vid_sram_raddr7 = vid_sram_raddr_total; vid_sram_raddr15 = vid_sram_raddr_total;
	end 
end 
always @* begin
	if(state == MASTER) begin
		n_interfinish =  interfinish | (tmpwaddr == 4'd15);
	end else begin 
		n_interfinish = 4'd0;
	end  
	if(state == MASTER) begin 
		if(tmpwaddr != 4'd15) n_tmpwaddr = tmpwaddr + 1;
		else n_tmpwaddr = tmpwaddr;
	end else begin 
		n_tmpwaddr = 4'd0;
	end 

	if(state == MASTER) begin
		if(interfinish == 0) begin 
			loc_sram_wen =  {K{1'b0}};
			loc_sram_waddr0 = tmpwaddr; 	loc_sram_wdata0 = 0;	loc_wbytemask0 = 0;
			loc_sram_waddr1 = tmpwaddr; 	loc_sram_wdata1 = 0;	loc_wbytemask1 = 0;
			loc_sram_waddr2 = tmpwaddr; 	loc_sram_wdata2 = 0;	loc_wbytemask2 = 0;
			loc_sram_waddr3 = tmpwaddr; 	loc_sram_wdata3 = 0;	loc_wbytemask3 = 0;
			loc_sram_waddr4 = tmpwaddr; 	loc_sram_wdata4 = 0;	loc_wbytemask4 = 0;
			loc_sram_waddr5 = tmpwaddr; 	loc_sram_wdata5 = 0;	loc_wbytemask5 = 0;
			loc_sram_waddr6 = tmpwaddr; 	loc_sram_wdata6 = 0;	loc_wbytemask6 = 0;
			loc_sram_waddr7 = tmpwaddr; 	loc_sram_wdata7 = 0;	loc_wbytemask7 = 0;
			loc_sram_waddr8 = tmpwaddr; 	loc_sram_wdata8 = 0;	loc_wbytemask8 = 0;
			loc_sram_waddr9 = tmpwaddr; 	loc_sram_wdata9 = 0;	loc_wbytemask9 = 0;
			loc_sram_waddr10 = tmpwaddr; 	loc_sram_wdata10 = 0;	loc_wbytemask10 = 0;
			loc_sram_waddr11 = tmpwaddr; 	loc_sram_wdata11 = 0;	loc_wbytemask11 = 0;
			loc_sram_waddr12 = tmpwaddr; 	loc_sram_wdata12 = 0;	loc_wbytemask12 = 0;
			loc_sram_waddr13 = tmpwaddr; 	loc_sram_wdata13 = 0;	loc_wbytemask13 = 0;
			loc_sram_waddr14 = tmpwaddr; 	loc_sram_wdata14 = 0;	loc_wbytemask14 = 0;
			loc_sram_waddr15 = tmpwaddr; 	loc_sram_wdata15 = 0;	loc_wbytemask15 = 0;
		end else begin
			loc_sram_wen = {K{master_locsram_wen}};
		 	loc_sram_waddr0 = master_loc_sram_waddr0; 		loc_sram_wdata0 = master_loc_sram_wdata0;	loc_wbytemask0 = master_loc_wbytemask0;
			loc_sram_waddr1 = master_loc_sram_waddr1; 		loc_sram_wdata1 = master_loc_sram_wdata1;	loc_wbytemask1 = master_loc_wbytemask1;
			loc_sram_waddr2 = master_loc_sram_waddr2; 		loc_sram_wdata2 = master_loc_sram_wdata2;	loc_wbytemask2 = master_loc_wbytemask2;
			loc_sram_waddr3 = master_loc_sram_waddr3; 		loc_sram_wdata3 = master_loc_sram_wdata3;	loc_wbytemask3 = master_loc_wbytemask3;
			loc_sram_waddr4 = master_loc_sram_waddr4; 		loc_sram_wdata4 = master_loc_sram_wdata4;	loc_wbytemask4 = master_loc_wbytemask4;
			loc_sram_waddr5 = master_loc_sram_waddr5; 		loc_sram_wdata5 = master_loc_sram_wdata5;	loc_wbytemask5 = master_loc_wbytemask5;
			loc_sram_waddr6 = master_loc_sram_waddr6; 		loc_sram_wdata6 = master_loc_sram_wdata6;	loc_wbytemask6 = master_loc_wbytemask6;
			loc_sram_waddr7 = master_loc_sram_waddr7; 		loc_sram_wdata7 = master_loc_sram_wdata7;	loc_wbytemask7 = master_loc_wbytemask7;
			loc_sram_waddr8 = master_loc_sram_waddr8; 		loc_sram_wdata8 = master_loc_sram_wdata8;	loc_wbytemask8 = master_loc_wbytemask8;
			loc_sram_waddr9 = master_loc_sram_waddr9; 		loc_sram_wdata9 = master_loc_sram_wdata9;	loc_wbytemask9 = master_loc_wbytemask9;
			loc_sram_waddr10 = master_loc_sram_waddr10; 	loc_sram_wdata10 = master_loc_sram_wdata10;	loc_wbytemask10 = master_loc_wbytemask10;
			loc_sram_waddr11 = master_loc_sram_waddr11; 	loc_sram_wdata11 = master_loc_sram_wdata11;	loc_wbytemask11 = master_loc_wbytemask11;
			loc_sram_waddr12 = master_loc_sram_waddr12; 	loc_sram_wdata12 = master_loc_sram_wdata12;	loc_wbytemask12 = master_loc_wbytemask12;
			loc_sram_waddr13 = master_loc_sram_waddr13; 	loc_sram_wdata13 = master_loc_sram_wdata13;	loc_wbytemask13 = master_loc_wbytemask13;
			loc_sram_waddr14 = master_loc_sram_waddr14; 	loc_sram_wdata14 = master_loc_sram_wdata14;	loc_wbytemask14 = master_loc_wbytemask14;
			loc_sram_waddr15 = master_loc_sram_waddr15; 	loc_sram_wdata15 = master_loc_sram_wdata15;	loc_wbytemask15 = master_loc_wbytemask15;
		end 
	end else begin 	
		loc_sram_wen =  {K{1'b1}};
		loc_sram_waddr0 = 0; 	loc_sram_wdata0 = 0;	loc_wbytemask0 = {D{1'b1}};
		loc_sram_waddr1 = 0; 	loc_sram_wdata1 = 0;	loc_wbytemask1 = {D{1'b1}};
		loc_sram_waddr2 = 0; 	loc_sram_wdata2 = 0;	loc_wbytemask2 = {D{1'b1}};
		loc_sram_waddr3 = 0; 	loc_sram_wdata3 = 0;	loc_wbytemask3 = {D{1'b1}};
		loc_sram_waddr4 = 0; 	loc_sram_wdata4 = 0;	loc_wbytemask4 = {D{1'b1}};
		loc_sram_waddr5 = 0; 	loc_sram_wdata5 = 0;	loc_wbytemask5 = {D{1'b1}};
		loc_sram_waddr6 = 0; 	loc_sram_wdata6 = 0;	loc_wbytemask6 = {D{1'b1}};
		loc_sram_waddr7 = 0; 	loc_sram_wdata7 = 0;	loc_wbytemask7 = {D{1'b1}};
		loc_sram_waddr8 = 0; 	loc_sram_wdata8 = 0;	loc_wbytemask8 = {D{1'b1}};
		loc_sram_waddr9 = 0; 	loc_sram_wdata9 = 0;	loc_wbytemask9 = {D{1'b1}};
		loc_sram_waddr10 = 0; 	loc_sram_wdata10 = 0;	loc_wbytemask10 = {D{1'b1}};
		loc_sram_waddr11 = 0; 	loc_sram_wdata11 = 0;	loc_wbytemask11 = {D{1'b1}};
		loc_sram_waddr12 = 0; 	loc_sram_wdata12 = 0;	loc_wbytemask12 = {D{1'b1}};
		loc_sram_waddr13 = 0; 	loc_sram_wdata13 = 0;	loc_wbytemask13 = {D{1'b1}};
		loc_sram_waddr14 = 0; 	loc_sram_wdata14 = 0;	loc_wbytemask14 = {D{1'b1}};
		loc_sram_waddr15 = 0; 	loc_sram_wdata15 = 0;	loc_wbytemask15 = {D{1'b1}};
	end 
end 

assign w0_vid_rdata = vid_sram_rdata0;
assign w1_vid_rdata = vid_sram_rdata1;
assign w2_vid_rdata = vid_sram_rdata2;
assign w3_vid_rdata = vid_sram_rdata3;
assign w4_vid_rdata = vid_sram_rdata4;
assign w5_vid_rdata = vid_sram_rdata5;
assign w6_vid_rdata = vid_sram_rdata6;
assign w7_vid_rdata = vid_sram_rdata7;
assign w8_vid_rdata = vid_sram_rdata8;
assign w9_vid_rdata = vid_sram_rdata9;
assign w10_vid_rdata = vid_sram_rdata10;
assign w11_vid_rdata = vid_sram_rdata11;
assign w12_vid_rdata = vid_sram_rdata12;
assign w13_vid_rdata = vid_sram_rdata13;
assign w14_vid_rdata = vid_sram_rdata14;
assign w15_vid_rdata = vid_sram_rdata15;

// dist sram write in
assign dist_sram_raddr0 = {vid0, sub_bat0};
assign dist_sram_raddr1 = {vid1, sub_bat1};
assign dist_sram_raddr2 = {vid2, sub_bat2};
assign dist_sram_raddr3 = {vid3, sub_bat3};
assign dist_sram_raddr4 = {vid4, sub_bat4};
assign dist_sram_raddr5 = {vid5, sub_bat5};
assign dist_sram_raddr6 = {vid6, sub_bat6};
assign dist_sram_raddr7 = {vid7, sub_bat7};
assign dist_sram_raddr8 = {vid8, sub_bat8};
assign dist_sram_raddr9 = {vid9, sub_bat9};
assign dist_sram_raddr10 = {vid10, sub_bat10};
assign dist_sram_raddr11 = {vid11, sub_bat11};
assign dist_sram_raddr12 = {vid12, sub_bat12};
assign dist_sram_raddr13 = {vid13, sub_bat13};
assign dist_sram_raddr14 = {vid14, sub_bat14};
assign dist_sram_raddr15 = {vid15, sub_bat15};

assign w0_dist_rdata = dist_sram_rdata0;
assign w1_dist_rdata = dist_sram_rdata1;
assign w2_dist_rdata = dist_sram_rdata2;
assign w3_dist_rdata = dist_sram_rdata3;
assign w4_dist_rdata = dist_sram_rdata4;
assign w5_dist_rdata = dist_sram_rdata5;
assign w6_dist_rdata = dist_sram_rdata6;
assign w7_dist_rdata = dist_sram_rdata7;
assign w8_dist_rdata = dist_sram_rdata8;
assign w9_dist_rdata = dist_sram_rdata9;
assign w10_dist_rdata = dist_sram_rdata10;
assign w11_dist_rdata = dist_sram_rdata11;
assign w12_dist_rdata = dist_sram_rdata12;
assign w13_dist_rdata = dist_sram_rdata13;
assign w14_dist_rdata = dist_sram_rdata14;
assign w15_dist_rdata = dist_sram_rdata15;


always@ (posedge clk) begin
	if (~rst_n) begin
		iter <= 4'd0;
		state <= IDLE;
		batch_num <= 8'd0;
		tmpwaddr <= 4'd0;
		interfinish <= 1'd0;
		part_finish <= 1'b0;
	end else begin
		iter <= n_iter;
		state <= n_state;
		batch_num <= n_batch_num;
		tmpwaddr <= n_tmpwaddr;
		interfinish <= n_interfinish;
		if(state == FIN) 
			part_finish <= 1;
	end
end

always@* begin 
	if(state == IDLE)  
		n_batch_num = batch_num;
	else  
		n_batch_num = (sub_bat0 == 4'd14) ? batch_num + 1 : batch_num;
end 

// FSM
always@* begin
	if(~rst_n) begin 
		rst_n_worker = 1'b0;
	end else begin 
		case(state) 
			IDLE: rst_n_worker = rst_n;
			WORKER: rst_n_worker = 1'b1;//batch_finish0 == 1 ? 1'b0 : 1'b1;
			MASTER: rst_n_worker = 1'b1;
			FIN: rst_n_worker = 1'b0;
		endcase 
	end 

	case(state)
		IDLE: begin
			en_worker = en;
			en_master = 0;
			//rst_n_worker = rst_n;
			rst_n_master = rst_n;
			if (en) begin
				n_state = WORKER;
			end else begin
				n_state = IDLE;
			end
			n_iter = iter;
		end
		WORKER: begin
			en_worker = en;
			en_master = 0;
			rst_n_master = 0;
			if (batch_finish0) begin
				n_state = MASTER;
				//rst_n_worker = 0;
			end else begin
				n_state = WORKER;
				//rst_n_worker = 1;
			end
			n_iter = iter;
		end
		MASTER: begin
			en_worker = 0;
			en_master = en && interfinish;
			//rst_n_worker = 0;
			if (master_finish) begin 
				n_state = FIN;
				rst_n_master = 0;
				n_iter = iter + 1;
			end else begin 
				n_state = MASTER; 
				rst_n_master = 1;
				n_iter = iter;
			end 
		end
		FIN: begin
			en_worker = 0;
			en_master = 0;
			//rst_n_worker = 0;
			rst_n_master = 0;
			n_state = IDLE;
			n_iter = iter;
		end
	endcase
end
endmodule 