module master_top #(
parameter Q = 16,
parameter PRO_BW = 8,
parameter NEXT_BW = 4,
parameter K = 16,
parameter VID_BW = 16,
parameter BUF_BW = 5, // log(2*Q)
parameter OFFSET_BW = 5, // 0-16 partial sum
parameter VID_ADDR_SPACE = 5,
parameter LOC_BW = 5,
parameter D = 256,
parameter LOC_ADDR_SPACE = 4
) (
input clk,
input rst_n, 
input enable,
// inputs 
input [NEXT_BW*Q-1:0] in_next_arr,
input [PRO_BW*K-1:0] in_mi_j, 
input [PRO_BW*K-1:0] in_mj_i, 
input [VID_BW*Q-1:0] in_v_gidx, 
input [PRO_BW*Q-1:0] in_proposal_nums,
// outputs 
output reg [7:0] epoch,
output reg [K-1:0] vidsram_wen, // 0 at MSB
output reg ready,
output reg finish,
// vidsram writing  
output [VID_BW*Q-1:0] vid_sram_wdata0,  output [VID_ADDR_SPACE-1:0] vid_sram_waddr0,
output [VID_BW*Q-1:0] vid_sram_wdata1,  output [VID_ADDR_SPACE-1:0] vid_sram_waddr1,
output [VID_BW*Q-1:0] vid_sram_wdata2,  output [VID_ADDR_SPACE-1:0] vid_sram_waddr2,
output [VID_BW*Q-1:0] vid_sram_wdata3,  output [VID_ADDR_SPACE-1:0] vid_sram_waddr3,
output [VID_BW*Q-1:0] vid_sram_wdata4,  output [VID_ADDR_SPACE-1:0] vid_sram_waddr4,
output [VID_BW*Q-1:0] vid_sram_wdata5,  output [VID_ADDR_SPACE-1:0] vid_sram_waddr5,
output [VID_BW*Q-1:0] vid_sram_wdata6,  output [VID_ADDR_SPACE-1:0] vid_sram_waddr6,
output [VID_BW*Q-1:0] vid_sram_wdata7,  output [VID_ADDR_SPACE-1:0] vid_sram_waddr7,
output [VID_BW*Q-1:0] vid_sram_wdata8,  output [VID_ADDR_SPACE-1:0] vid_sram_waddr8,
output [VID_BW*Q-1:0] vid_sram_wdata9,  output [VID_ADDR_SPACE-1:0] vid_sram_waddr9,
output [VID_BW*Q-1:0] vid_sram_wdata10, output [VID_ADDR_SPACE-1:0] vid_sram_waddr10,
output [VID_BW*Q-1:0] vid_sram_wdata11, output [VID_ADDR_SPACE-1:0] vid_sram_waddr11,
output [VID_BW*Q-1:0] vid_sram_wdata12, output [VID_ADDR_SPACE-1:0] vid_sram_waddr12,
output [VID_BW*Q-1:0] vid_sram_wdata13, output [VID_ADDR_SPACE-1:0] vid_sram_waddr13,
output [VID_BW*Q-1:0] vid_sram_wdata14, output [VID_ADDR_SPACE-1:0] vid_sram_waddr14,
output [VID_BW*Q-1:0] vid_sram_wdata15, output [VID_ADDR_SPACE-1:0] vid_sram_waddr15
// loc sram writing 

);
wire pingpong = 0;
localparam IDLE=2'd0, RUNS=2'd1, DELAY=2'd2, FINISH=2'd3;
localparam PSUM_READY = 3;
localparam DONEII = 6;
reg [1:0] nstate, state;
// reg rst_n, enable;
// localparam WDATII = 6; // WDATII = PSUM_READY + 3
// epoch[7:4] -> i, current partition
reg [2:0] delay, n_delay;
reg [7:0] n_epoch;
reg [NEXT_BW-1:0] next_arr[0:Q-1];      // register             
reg [PRO_BW-1:0] proposal_nums[0:Q-1];  // register         
reg [PRO_BW-1:0] mi_j[0:K-1];           // register 
reg [PRO_BW-1:0] mj_i[0:K-1];           // register 
reg [NEXT_BW-1:0] real_next_arr[0:Q-1], nreal_next_arr[0:Q-1], buff_1_next[0:Q-1], buff_next[0:Q-1];

// vid sram
reg [Q*VID_BW-1:0] vidsram_wdata[0:K-1];
reg [VID_ADDR_SPACE-1:0] vidsram_waddr[0:K-1];
// loc sram
reg [D*LOC_BW-1:0] locsram_wdata[0:Q-1];
reg locsram_wen[0:Q-1];
reg [D-1:0] locsram_wbytemask[0:Q-1], n_locsram_wbytemask[0:Q-1];
reg [LOC_ADDR_SPACE-1:0] locsram_addr[0:Q-1];

// sram wire connect
assign vid_sram_wdata0 = vidsram_wdata[0];    assign vid_sram_waddr0 =   vidsram_waddr[0];   
assign vid_sram_wdata1 = vidsram_wdata[1];    assign vid_sram_waddr1 =   vidsram_waddr[1];   
assign vid_sram_wdata2 = vidsram_wdata[2];    assign vid_sram_waddr2 =   vidsram_waddr[2];   
assign vid_sram_wdata3 = vidsram_wdata[3];    assign vid_sram_waddr3 =   vidsram_waddr[3];   
assign vid_sram_wdata4 = vidsram_wdata[4];    assign vid_sram_waddr4 =   vidsram_waddr[4];   
assign vid_sram_wdata5 = vidsram_wdata[5];    assign vid_sram_waddr5 =   vidsram_waddr[5];   
assign vid_sram_wdata6 = vidsram_wdata[6];    assign vid_sram_waddr6 =   vidsram_waddr[6];   
assign vid_sram_wdata7 = vidsram_wdata[7];    assign vid_sram_waddr7 =   vidsram_waddr[7];   
assign vid_sram_wdata8 = vidsram_wdata[8];    assign vid_sram_waddr8 =   vidsram_waddr[8];   
assign vid_sram_wdata9 = vidsram_wdata[9];    assign vid_sram_waddr9 =   vidsram_waddr[9];   
assign vid_sram_wdata10 = vidsram_wdata[10];  assign vid_sram_waddr10 =  vidsram_waddr[10];       
assign vid_sram_wdata11 = vidsram_wdata[11];  assign vid_sram_waddr11 =  vidsram_waddr[11];       
assign vid_sram_wdata12 = vidsram_wdata[12];  assign vid_sram_waddr12 =  vidsram_waddr[12];       
assign vid_sram_wdata13 = vidsram_wdata[13];  assign vid_sram_waddr13 =  vidsram_waddr[13];       
assign vid_sram_wdata14 = vidsram_wdata[14];  assign vid_sram_waddr14 =  vidsram_waddr[14];       
assign vid_sram_wdata15 = vidsram_wdata[15];  assign vid_sram_waddr15 =  vidsram_waddr[15];       
// ================================================
// TOOD: prepare: next_arr, mi_j, mj_i, v_gidx , proposal_nums

// ================================================
reg [VID_BW-1:0] v_gidx[0:Q-1]; // registers, from vid sram
// K buffers, each of Q 
reg [VID_BW-1:0] buffer [0:K-1] [0:2*Q-1], n_buffer[0:K-1][0:2*Q-1];
reg [BUF_BW-1:0] accum[0:K-1], n_accum[0:K-1]; // buffer size for each of K buffers
reg [BUF_BW-1:0] buffer_idx[0:Q-1], nbuffer_idx[0:Q-1]; // additioanl bit??
reg export[0:K-1], n_export[0:K-1];
reg [BUF_BW-1:0] buffaccum[0:K-1], n_buffaccum[0:K-1]; // for buffer indexing's accum
reg [K-1:0] onehot[0:Q-1];
reg [OFFSET_BW-1:0] partial_sum[0:Q-1][0:K-1],n_partial_sum[0:Q-1][0:K-1];
reg psum_set, n_psum_set;
integer o_idx, in_idx;
integer accumidx;
integer partial_i, partial_j, check_i;
integer buffi,buffj;

always @* begin 
    if(~enable) n_psum_set = 0;
    else begin 
        if(state == RUNS && epoch == PSUM_READY) n_psum_set = 1;
        else n_psum_set = psum_set;
    end 
    if(~enable) n_delay = 0;
    else begin 
        if(state == DELAY)  n_delay = delay + 1;
        else                n_delay = delay;
    end 
    if(~enable) n_epoch = 0;
    else begin 
        if(state == RUNS && epoch < 8'd255) n_epoch = epoch + 1;
        else              n_epoch = epoch; 
    end 

    for(o_idx = 0; o_idx < Q; o_idx = o_idx + 1) begin 
        for(in_idx = 0; in_idx < K; in_idx = in_idx + 1) begin
            onehot[o_idx][in_idx] = real_next_arr[o_idx] == in_idx;
        end 
    end 
    
    for(partial_j = 0; partial_j < K; partial_j = partial_j + 1) begin
        n_partial_sum[0][partial_j] =  onehot[0][partial_j];
        n_partial_sum[1][partial_j] =  onehot[0][partial_j]+onehot[1][partial_j];
        n_partial_sum[2][partial_j] =  onehot[0][partial_j]+onehot[1][partial_j]+onehot[2][partial_j];
        n_partial_sum[3][partial_j] =  onehot[0][partial_j]+onehot[1][partial_j]+onehot[2][partial_j]+onehot[3][partial_j];
        n_partial_sum[4][partial_j] =  onehot[0][partial_j]+onehot[1][partial_j]+onehot[2][partial_j]+onehot[3][partial_j]+onehot[4][partial_j];
        n_partial_sum[5][partial_j] =  onehot[0][partial_j]+onehot[1][partial_j]+onehot[2][partial_j]+onehot[3][partial_j]+onehot[4][partial_j]+onehot[5][partial_j];
        n_partial_sum[6][partial_j] =  onehot[0][partial_j]+onehot[1][partial_j]+onehot[2][partial_j]+onehot[3][partial_j]+onehot[4][partial_j]+onehot[5][partial_j]+onehot[6][partial_j];
        n_partial_sum[7][partial_j] =  onehot[0][partial_j]+onehot[1][partial_j]+onehot[2][partial_j]+onehot[3][partial_j]+onehot[4][partial_j]+onehot[5][partial_j]+onehot[6][partial_j]+onehot[7][partial_j];
        n_partial_sum[8][partial_j] =  onehot[0][partial_j]+onehot[1][partial_j]+onehot[2][partial_j]+onehot[3][partial_j]+onehot[4][partial_j]+onehot[5][partial_j]+onehot[6][partial_j]+onehot[7][partial_j]+onehot[8][partial_j];
        n_partial_sum[9][partial_j] =  onehot[0][partial_j]+onehot[1][partial_j]+onehot[2][partial_j]+onehot[3][partial_j]+onehot[4][partial_j]+onehot[5][partial_j]+onehot[6][partial_j]+onehot[7][partial_j]+onehot[8][partial_j]+onehot[9][partial_j];
        n_partial_sum[10][partial_j] = onehot[0][partial_j]+onehot[1][partial_j]+onehot[2][partial_j]+onehot[3][partial_j]+onehot[4][partial_j]+onehot[5][partial_j]+onehot[6][partial_j]+onehot[7][partial_j]+onehot[8][partial_j]+onehot[9][partial_j]+onehot[10][partial_j];
        n_partial_sum[11][partial_j] = onehot[0][partial_j]+onehot[1][partial_j]+onehot[2][partial_j]+onehot[3][partial_j]+onehot[4][partial_j]+onehot[5][partial_j]+onehot[6][partial_j]+onehot[7][partial_j]+onehot[8][partial_j]+onehot[9][partial_j]+onehot[10][partial_j]+onehot[11][partial_j];
        n_partial_sum[12][partial_j] = onehot[0][partial_j]+onehot[1][partial_j]+onehot[2][partial_j]+onehot[3][partial_j]+onehot[4][partial_j]+onehot[5][partial_j]+onehot[6][partial_j]+onehot[7][partial_j]+onehot[8][partial_j]+onehot[9][partial_j]+onehot[10][partial_j]+onehot[11][partial_j]+onehot[12][partial_j];
        n_partial_sum[13][partial_j] = onehot[0][partial_j]+onehot[1][partial_j]+onehot[2][partial_j]+onehot[3][partial_j]+onehot[4][partial_j]+onehot[5][partial_j]+onehot[6][partial_j]+onehot[7][partial_j]+onehot[8][partial_j]+onehot[9][partial_j]+onehot[10][partial_j]+onehot[11][partial_j]+onehot[12][partial_j]+onehot[13][partial_j];
        n_partial_sum[14][partial_j] = onehot[0][partial_j]+onehot[1][partial_j]+onehot[2][partial_j]+onehot[3][partial_j]+onehot[4][partial_j]+onehot[5][partial_j]+onehot[6][partial_j]+onehot[7][partial_j]+onehot[8][partial_j]+onehot[9][partial_j]+onehot[10][partial_j]+onehot[11][partial_j]+onehot[12][partial_j]+onehot[13][partial_j]+onehot[14][partial_j];
        n_partial_sum[15][partial_j] = onehot[0][partial_j]+onehot[1][partial_j]+onehot[2][partial_j]+onehot[3][partial_j]+onehot[4][partial_j]+onehot[5][partial_j]+onehot[6][partial_j]+onehot[7][partial_j]+onehot[8][partial_j]+onehot[9][partial_j]+onehot[10][partial_j]+onehot[11][partial_j]+onehot[12][partial_j]+onehot[13][partial_j]+onehot[14][partial_j]+onehot[15][partial_j];
    
    end 
    // ----------- same time to write into ----------------
    for(partial_i = 0; partial_i < Q; partial_i = partial_i + 1) begin
        if(psum_set) 
        nbuffer_idx[partial_i] = (partial_sum[partial_i][buff_1_next[partial_i]] - 1) + (accum[buff_1_next[partial_i]] >= Q ? accum[buff_1_next[partial_i]] - Q : accum[buff_1_next[partial_i]]) ;
        else 
        nbuffer_idx[partial_i] = buffer_idx[partial_i];
        // TODO: accum[q] == Q also update to partial_sum[15][q], / transfer out 
    end
       
    for(accumidx = 0; accumidx < K; accumidx = accumidx + 1) begin 
        n_buffaccum[accumidx] = accum[accumidx] >= Q ? accum[accumidx] - Q : accum[accumidx]; // retain the offset that to be FIFOed

        if(psum_set) begin 
            if(accum[accumidx] >= Q) begin 
                n_accum[accumidx] = accum[accumidx] - Q + partial_sum[Q-1][accumidx]; // partial sum !!!! ;// check_acc[accumidx] - Q;
                n_export[accumidx] = 1;
            end else begin 
                n_accum[accumidx] = accum[accumidx] + partial_sum[Q-1][accumidx];//accum[accumidx];//check_acc[accumidx];
                n_export[accumidx] = 0;
            end
        end else begin 
            n_export[accumidx] = export[accumidx];
            n_accum[accumidx] = accum[accumidx];
        end  
    
    end 
    // -------------------------------------------
    for(buffi = 0; buffi < K; buffi = buffi + 1) begin 
        for(buffj = 0; buffj < 2*Q; buffj = buffj + 1) begin  
            if(psum_set) begin 
                if(buffj < Q && export[buffi] == 1 && buffj < buffaccum[buffi]) begin 
                    // shift 
                    n_buffer[buffi][buffj] = buffer[buffi][buffj + Q];
                end else begin 
                    // take new 
                    if(buffj < buffaccum[buffi]) begin
                        n_buffer[buffi][buffj] = buffer[buffi][buffj]; 
                    end else begin 
                        n_buffer[buffi][buffj] =
                                            ((buff_next[0] == buffi) * (buffer_idx[0] == buffj) * v_gidx[0]) |
                                            ((buff_next[1] == buffi) * (buffer_idx[1] == buffj) * v_gidx[1]) |
                                            ((buff_next[2] == buffi) * (buffer_idx[2] == buffj) * v_gidx[2]) |
                                            ((buff_next[3] == buffi) * (buffer_idx[3] == buffj) * v_gidx[3]) |
                                            ((buff_next[4] == buffi) * (buffer_idx[4] == buffj) * v_gidx[4]) |
                                            ((buff_next[5] == buffi) * (buffer_idx[5] == buffj) * v_gidx[5]) |
                                            ((buff_next[6] == buffi) * (buffer_idx[6] == buffj) * v_gidx[6]) |
                                            ((buff_next[7] == buffi) * (buffer_idx[7] == buffj) * v_gidx[7]) |
                                            ((buff_next[8] == buffi) * (buffer_idx[8] == buffj) * v_gidx[8]) |
                                            ((buff_next[9] == buffi) * (buffer_idx[9] == buffj) * v_gidx[9]) |
                                            ((buff_next[10] == buffi) * (buffer_idx[10] == buffj) * v_gidx[10]) |
                                            ((buff_next[11] == buffi) * (buffer_idx[11] == buffj) * v_gidx[11]) |
                                            ((buff_next[12] == buffi) * (buffer_idx[12] == buffj) * v_gidx[12]) |
                                            ((buff_next[13] == buffi) * (buffer_idx[13] == buffj) * v_gidx[13]) |
                                            ((buff_next[14] == buffi) * (buffer_idx[14] == buffj) * v_gidx[14]) |
                                            ((buff_next[15] == buffi) * (buffer_idx[15] == buffj) * v_gidx[15]);
                    end 
                end 
            end else begin 
                n_buffer[buffi][buffj] = buffer[buffi][buffj];
            end 
        end 
    end 

end 

// comb7 get xij
reg [PRO_BW-1:0] xijs[0:K-1]; // n_xijs[0:K-1];

integer j, qiter;
wire [7:0] tmpepoch = epoch >= 2 ? epoch - 2 : epoch;
always @* begin 
    for(j = 0; j < K; j = j + 1) begin 
        xijs[j] = mi_j[j] < mj_i[j] ? mi_j[j] : mj_i[j];
    end 
    for(qiter = 0; qiter < Q; qiter = qiter + 1) begin
        nreal_next_arr[qiter] = xijs[next_arr[qiter]] > proposal_nums[qiter] ? next_arr[qiter] : tmpepoch[7:4]; // < xij move, if not stay at current 
    end 
end 
integer mask_i;
always @* begin 
    for(mask_i = 0; mask_i < Q; mask_i = mask_i + 1) begin 
        (* synthesis, parallel_case *)
        case(v_gidx[mask_i][7:0])
            0:    n_locsram_wbytemask[mask_i] = 256'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            1:    n_locsram_wbytemask[mask_i] = 256'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            2:    n_locsram_wbytemask[mask_i] = 256'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            3:    n_locsram_wbytemask[mask_i] = 256'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            4:    n_locsram_wbytemask[mask_i] = 256'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            5:    n_locsram_wbytemask[mask_i] = 256'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            6:    n_locsram_wbytemask[mask_i] = 256'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            7:    n_locsram_wbytemask[mask_i] = 256'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            8:    n_locsram_wbytemask[mask_i] = 256'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            9:    n_locsram_wbytemask[mask_i] = 256'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            10:   n_locsram_wbytemask[mask_i] = 256'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            11:   n_locsram_wbytemask[mask_i] = 256'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            12:   n_locsram_wbytemask[mask_i] = 256'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            13:   n_locsram_wbytemask[mask_i] = 256'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            14:   n_locsram_wbytemask[mask_i] = 256'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            15:   n_locsram_wbytemask[mask_i] = 256'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            16:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            17:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            18:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            19:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            20:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            21:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            22:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            23:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            24:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            25:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            26:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            27:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            28:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            29:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            30:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            31:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            33:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            34:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            35:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            36:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            37:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            38:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            39:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            40:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            41:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            42:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            43:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            44:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            45:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            46:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            47:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            48:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            49:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            50:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            51:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            52:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            53:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            54:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            55:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            56:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            57:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            58:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            59:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            60:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            61:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            62:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            63:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            64:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            65:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            66:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            67:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            68:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            69:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            70:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            71:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            72:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            73:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            74:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            75:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            76:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            77:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            78:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            79:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            80:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            81:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            82:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            83:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            84:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            85:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            86:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            87:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            88:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            89:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            90:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            91:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            92:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            93:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            94:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            95:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            96:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            97:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            98:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            99:   n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            100:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            101:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            102:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            103:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            104:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            105:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            106:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            107:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            108:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            109:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            110:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            111:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            112:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            113:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            114:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            115:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            116:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            117:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            118:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            119:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            120:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            121:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            122:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            123:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            124:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            125:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            126:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            127:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            128:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            129:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            130:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            131:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            132:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            133:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            134:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            135:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            136:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            137:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            138:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            139:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            140:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            141:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            142:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            143:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            144:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            145:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            146:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            147:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            148:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            149:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            150:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            151:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            152:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            153:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            154:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            155:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            156:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            157:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            158:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            159:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            160:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            161:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            162:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            163:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            164:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            165:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            166:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            167:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            168:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            169:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            170:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            171:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            172:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            173:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            174:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            175:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
            176:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000;
            177:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000;
            178:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000;
            179:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000;
            180:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000;
            181:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;
            182:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000;
            183:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
            184:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000;
            185:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000;
            186:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000;
            187:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000;
            188:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000;
            189:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000;
            190:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000;
            191:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000;
            192:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000;
            193:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000;
            194:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000;
            195:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000;
            196:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000;
            197:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000;
            198:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000;
            199:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000;
            200:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000;
            201:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000;
            202:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000;
            203:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000;
            204:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000;
            205:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000;
            206:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000;
            207:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000;
            208:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000;
            209:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000;
            210:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000;
            211:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000;
            212:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000;
            213:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000;
            214:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000;
            215:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
            216:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000;
            217:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000;
            218:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000;
            219:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000;
            220:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000;
            221:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000;
            222:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000;
            223:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000;
            224:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000;
            225:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000;
            226:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000;
            227:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000;
            228:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000;
            229:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000;
            230:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000;
            231:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000;
            232:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000;
            233:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000;
            234:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000;
            235:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000;
            236:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000;
            237:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000;
            238:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000;
            239:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000;
            240:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000;
            241:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000;
            242:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000;
            243:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000;
            244:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000;
            245:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000;
            246:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000;
            247:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000;
            248:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000;
            249:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000;
            250:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000;
            251:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
            252:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
            253:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100;
            254:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;
            255:  n_locsram_wbytemask[mask_i] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
        endcase 
    end 
end 
// total epoch = N(4096) / Q(16)
integer loci;
integer export_i;
integer ri, rk, rj, si, sk, sq, pi, pj;
always @* begin 
    if(~enable) begin 
        nstate = IDLE;
    end else begin 
        case(state) 
            IDLE: nstate = RUNS;
            RUNS: nstate = (epoch == 8'd255) ? DELAY : RUNS;
            DELAY: nstate = (delay == DONEII) ? FINISH : DELAY;
            FINISH: nstate = FINISH;
        endcase 
    end 
end 
always @(posedge clk) begin 
    if(~rst_n) begin 
        state <= IDLE;
        psum_set <= 0;
        for(ri = 0; ri < Q; ri = ri + 1) begin 
            next_arr[ri] <= {NEXT_BW{1'b0}};
            proposal_nums[ri] <= {PRO_BW{1'b0}};
            v_gidx[ri] <= {VID_BW{1'b0}};
            real_next_arr[ri] <= {NEXT_BW{1'b0}};
            buff_next[ri] <= {NEXT_BW{1'b0}};
            buff_1_next[ri] <= {NEXT_BW{1'b0}};
            for(rj = 0; rj < K; rj = rj + 1) begin 
                buffer[rj][2*ri] <= {VID_BW{1'b0}};
                buffer[rj][2*ri+1] <= {VID_BW{1'b0}};
                partial_sum[ri][rj] <= {OFFSET_BW{1'b0}};
            end 
            buffer_idx[ri] <= {BUF_BW{1'b0}};
        end 
        vidsram_wen <= {K{1'b1}};
        for(rk = 0; rk < K; rk = rk + 1) begin 
            mi_j[rk] <= {PRO_BW{1'b0}};
            mj_i[rk] <= {PRO_BW{1'b0}};
            vidsram_wdata[rk] <= {Q*VID_BW-1{1'b0}};
            vidsram_waddr[rk] <= {VID_ADDR_SPACE{1'b0}};
            accum[rk] <= {BUF_BW{1'b0}};
            export[rk] <= 1'b0;
            buffaccum[rk] <= {BUF_BW{1'b0}};
        end 
        epoch <= 0;
        ready <= 0;
        finish <= 0;
        delay <= 0;
    end else begin
        state <= nstate; 
        epoch <= n_epoch;
        // $write("epoch: %d\n",epoch);
        delay <= n_delay;
        psum_set <= n_psum_set;
        if(state == FINISH) finish <= 1;
        else                finish <= 0;
        {next_arr[0],next_arr[1],next_arr[2],next_arr[3],next_arr[4],next_arr[5],next_arr[6],next_arr[7],
        next_arr[8],next_arr[9],next_arr[10],next_arr[11],next_arr[12],next_arr[13],next_arr[14],next_arr[15]}
            <= in_next_arr;
        {proposal_nums[0],proposal_nums[1],proposal_nums[2],proposal_nums[3],proposal_nums[4],proposal_nums[5],proposal_nums[6],proposal_nums[7],
        proposal_nums[8],proposal_nums[9],proposal_nums[10],proposal_nums[11],proposal_nums[12],proposal_nums[13],proposal_nums[14],proposal_nums[15]}
            <= in_proposal_nums;
        {v_gidx[0],v_gidx[1],v_gidx[2],v_gidx[3],v_gidx[4],v_gidx[5],v_gidx[6],v_gidx[7],
        v_gidx[8],v_gidx[9],v_gidx[10],v_gidx[11],v_gidx[12],v_gidx[13],v_gidx[14],v_gidx[15]} 
            <= in_v_gidx;
        for(si = 0; si < Q; si = si + 1) begin 
            real_next_arr[si] <= nreal_next_arr[si];
            buff_1_next[si]<= real_next_arr[si];
            buff_next[si] <= buff_1_next[si];
            buffer_idx[si] <= nbuffer_idx[si];
        end 
        for(pi = 0; pi < Q; pi = pi + 1) begin 
            for(pj = 0; pj < K; pj = pj + 1) begin
                 partial_sum[pi][pj] <= n_partial_sum[pi][pj];
            end 
        end 

        {mi_j[0],mi_j[1],mi_j[2],mi_j[3],mi_j[4],mi_j[5],mi_j[6],mi_j[7],
        mi_j[8],mi_j[9],mi_j[10],mi_j[11],mi_j[12],mi_j[13],mi_j[14],mi_j[15]} <= in_mi_j;
        {mj_i[0],mj_i[1],mj_i[2],mj_i[3],mj_i[4],mj_i[5],mj_i[6],mj_i[7],
        mj_i[8],mj_i[9],mj_i[10],mj_i[11],mj_i[12],mj_i[13],mj_i[14],mj_i[15]} <= in_mj_i;
        if(enable && epoch > 4)
            ready <= 1;
        else 
            ready <= 0;
        for(sk = 0; sk < K; sk = sk + 1) begin 
            if(~enable) begin
                accum[sk] <= {BUF_BW{1'b0}};
                export[sk] <= 1'b0;
                buffaccum[sk] <= {BUF_BW{1'b0}};
            end else begin 
                accum[sk] <= n_accum[sk];
                export[sk] <= n_export[sk];
                buffaccum[sk] <= n_buffaccum[sk];
            end 
            for(sq = 0; sq < 2*Q; sq = sq + 1) begin 
                if(~enable) buffer[sk][sq] <= 0;
                else buffer[sk][sq] <= n_buffer[sk][sq];
            end 
        end 

        // write vid sram 
        for(export_i = 0; export_i < K; export_i = export_i + 1) begin 
            if(enable && state >= RUNS) begin 
                if(vidsram_wen[export_i] == 1'b0)  
                    vidsram_waddr[export_i]  <= vidsram_waddr[export_i] + 1;
                if(export[export_i] == 1) begin 
                    vidsram_wdata[export_i]  <= {buffer[export_i][0],buffer[export_i][1],buffer[export_i][2],buffer[export_i][3],buffer[export_i][4],buffer[export_i][5],buffer[export_i][6],buffer[export_i][7],buffer[export_i][8],buffer[export_i][9],buffer[export_i][10],buffer[export_i][11],buffer[export_i][12],buffer[export_i][13],buffer[export_i][14],buffer[export_i][15]};
                    vidsram_wen[export_i]  <= 1'b0;
                end else begin 
                    vidsram_wen[export_i]  <= 1'b1;
                end 
            end else begin 
                vidsram_wen[export_i]  <= 1'b1;
                vidsram_waddr[export_i] <= 5'd16 & {5{pingpong}};
            end 
            // if(vidsram_wen[export_i] !== 0) begin 
            //     $write(":epoch %d exportout target %d wen %h wdata %h\n", epoch, export_i, vidsram_wen[export_i], vidsram_wdata[export_i]);
            // end 
        end 
    
    

        // write loc sram
        if(epoch > 3) begin 
            // next_arr -> next_real_arr -> buff_next 
            for(loci = 0; loci < Q; loci = loci + 1) begin 
                locsram_wdata[loci] <= {D{1'b1, buff_next[loci]}};
                locsram_wbytemask[loci] <= n_locsram_wbytemask[loci];
                locsram_wen[loci] <= 1;
                // locsram_addr[loci] <= v_gidx[mask_i][D+3:D];  // TO MODIFIED
            end
            // TODO: start update read_waddr of vid ! 
        end

    end 
end 


endmodule





// case(next_arr[o_idx])
//     4'd0: onehot[o_idx] = 16'b0000000000000001;
//     4'd1: onehot[o_idx] = 16'b0000000000000010;
//     4'd2: onehot[o_idx] = 16'b0000000000000100;
// endcase 