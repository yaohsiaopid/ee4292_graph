module worker
#(
    parameter K = 16,
    parameter D = 256,
    parameter DIST_BW = 1,
    parameter DIST_ADDR_SPACE = 16,
    parameter LOC_BW = 5,
    parameter LOC_ADDR_SPACE = 4,
    parameter NEXT_BW = 4,
    parameter NEXT_ADDR_SPACE = 4,
    parameter PRO_BW = 8,
    parameter PRO_ADDR_SPACE = 4,
    parameter VID_BW = 16,  // 12???
    parameter VID_ADDR_SPACE = 4,
    parameter Q = 16,
	parameter WORK_IDX = 0
)
(
    input clk,
    input en,
    input rst_n,
    input [7:0] batch_num,
    input [Q*VID_BW-1:0] vid_rdata,					// 256
    input [D*DIST_BW-1:0] dist_rdata,				// 256
    input [D*(LOC_BW-1)-1:0] loc_rdata,             // input 256 X 4bit valid locations selected from top module

	output reg [3:0] sub_bat,						// 4
    output reg [VID_BW-1:0] vid,					// 16
	output reg [Q-1:0] next_bytemask,				// 16
    output reg [Q*NEXT_BW-1:0] next_wdata,			// 64
    output reg [NEXT_ADDR_SPACE-1:0] next_waddr,	// 4
	output reg [Q-1:0] pro_bytemask,				// 16
    output reg [Q*PRO_BW-1:0] pro_wdata,			// 128
	output reg [PRO_ADDR_SPACE-1:0] pro_waddr,		//4
    output reg ready,       // for part_reg[0:K-1]	// 1
    output reg batch_finish, // for next / proposal number	// 1
	output reg wen									// 1
);

// reg [15:0] vid;
reg [7:0] batch_num_reg;
reg [3:0] n_sub_bat;

reg [VID_BW-1:0] vid_reg [0:Q-1];
reg [VID_BW-1:0] n_vid;

reg [D-1:0] dist_reg;

reg [LOC_BW-2:0] loc_reg [0:D-1];

reg [K-1:0] n_loc_oh_reg [0:D-1];
reg [K-1:0] loc_oh_reg [0:D-1];

reg [4:0] dsum_reg [0:8*K-1];       // 256 / 32 = 8
reg [4:0] n_dsum_reg [0:8*K-1];       // 256 / 32 = 8

reg [7:0] part_reg [0:K-1];
reg [7:0] n_part_reg [0:K-1];

reg [Q*NEXT_BW-1:0] n_next_wdata;
reg [Q-1:0] n_next_bytemask;
reg [NEXT_ADDR_SPACE-1:0] n_next_waddr;

reg [Q*PRO_BW-1:0] n_pro_wdata;
reg [PRO_ADDR_SPACE-1:0] n_pro_waddr;
reg [Q-1:0] n_pro_bytemask;

reg [2:0] state, n_state;
reg n_batch_finish, n_ready;

reg [11:0] res0_comp [0:7];
reg [11:0] res1_comp [0:3];
reg [11:0] res2_comp [0:1];
reg [11:0] res3_comp;
reg [3:0] res4_comp;

reg [7:0] n_proposal_cnt [0:15];
reg [7:0] proposal_cnt [0:15];

reg part_en;

reg rst_n_in, en_in, n_wen;

integer i;

parameter IDLE = 3'd0, DELAY1 = 3'd1, SUB = 3'd2, DELAY2 = 3'd3, CHECK = 3'd4, FIN = 3'd5;

// batch_num, sub_bat, state, controls
always@(posedge clk) begin
	rst_n_in <= rst_n;
    if(~rst_n) begin
        next_wdata <= 64'd0;
        next_waddr <= 4'd0;
		next_bytemask <= 16'b1111_1111_1111_1111;
        pro_waddr <= 4'd0;
        pro_wdata <= 128'd0;
		pro_bytemask <= 16'b1111_1111_1111_1111;
        batch_num_reg <= 8'd0;
        sub_bat <= 4'd0;
        state <= 2'd0;
        batch_finish <= 1'd0;
        ready <= 1'd0;
		part_en <= 1'b0;
		res4_comp <= 4'd0;
		wen <= 1'd0;
		en_in <= 1'd0;
    end else begin
        next_waddr <= n_next_waddr;
		next_bytemask <= n_next_bytemask;
        next_wdata <= n_next_wdata;
		pro_waddr <= n_pro_waddr;
        pro_wdata <= n_pro_wdata;
		pro_bytemask <= n_pro_bytemask;
        batch_num_reg <= batch_num;
        sub_bat <= n_sub_bat;
        state <= n_state;
        batch_finish <= n_batch_finish;
        ready <= n_ready;
		part_en <= (batch_num_reg == 0 && sub_bat == 2) ? 1 : ready;
		res4_comp <= (res3_comp[11:4] > part_reg[WORK_IDX]) ? res3_comp[3:0] : WORK_IDX;
		wen <= n_wen;
		en_in <= en;
    end
end

// vid_reg, vid
always@(posedge clk) begin
	if(state == IDLE) begin
	    {vid_reg[0], vid_reg[1], vid_reg[2], vid_reg[3]} <= {vid_rdata[255:240], vid_rdata[239:224], vid_rdata[223:208], vid_rdata[207:192]};
        {vid_reg[4], vid_reg[5], vid_reg[6], vid_reg[7]} <= {vid_rdata[191:176], vid_rdata[175:160], vid_rdata[159:144], vid_rdata[143:128]};
        {vid_reg[8], vid_reg[9], vid_reg[10], vid_reg[11]} <= {vid_rdata[127:112], vid_rdata[111:96], vid_rdata[95:80], vid_rdata[79:64]};
        {vid_reg[12], vid_reg[13], vid_reg[14], vid_reg[15]} <= {vid_rdata[63:48], vid_rdata[47:32], vid_rdata[31:16], vid_rdata[15:0]};
        vid <= n_vid;
    end else if(batch_num_reg[3:0] != 4'b1111) begin
        {vid_reg[0], vid_reg[1], vid_reg[2], vid_reg[3]} <= {vid_reg[0], vid_reg[1], vid_reg[2], vid_reg[3]};
        {vid_reg[4], vid_reg[5], vid_reg[6], vid_reg[7]} <= {vid_reg[4], vid_reg[5], vid_reg[6], vid_reg[7]};
        {vid_reg[8], vid_reg[9], vid_reg[10], vid_reg[11]} <= {vid_reg[8], vid_reg[9], vid_reg[10], vid_reg[11]};
        {vid_reg[12], vid_reg[13], vid_reg[14], vid_reg[15]} <= {vid_reg[12], vid_reg[13], vid_reg[14], vid_reg[15]};
        vid <= n_vid;
    end else begin
        if(~rst_n_in) begin
            {vid_reg[0], vid_reg[1], vid_reg[2], vid_reg[3]} <= {16'd0, 16'd0, 16'd0, 16'd0};
            {vid_reg[4], vid_reg[5], vid_reg[6], vid_reg[7]} <= {16'd0, 16'd0, 16'd0, 16'd0};
            {vid_reg[8], vid_reg[9], vid_reg[10], vid_reg[11]} <= {16'd0, 16'd0, 16'd0, 16'd0};
            {vid_reg[12], vid_reg[13], vid_reg[14], vid_reg[15]} <= {16'd0, 16'd0, 16'd0, 16'd0};
            vid <= 16'd0;
        end else begin
            {vid_reg[0], vid_reg[1], vid_reg[2], vid_reg[3]} <= {vid_rdata[255:240], vid_rdata[239:224], vid_rdata[223:208], vid_rdata[207:192]};
            {vid_reg[4], vid_reg[5], vid_reg[6], vid_reg[7]} <= {vid_rdata[191:176], vid_rdata[175:160], vid_rdata[159:144], vid_rdata[143:128]};
            {vid_reg[8], vid_reg[9], vid_reg[10], vid_reg[11]} <= {vid_rdata[127:112], vid_rdata[111:96], vid_rdata[95:80], vid_rdata[79:64]};
            {vid_reg[12], vid_reg[13], vid_reg[14], vid_reg[15]} <= {vid_rdata[63:48], vid_rdata[47:32], vid_rdata[31:16], vid_rdata[15:0]};
            vid <= n_vid;
        end
    end
end

always@(posedge clk) begin
	if(~rst_n_in) begin
		for(i = 0; i < 16; i = i + 1) begin
			proposal_cnt[i] <= 8'd0;
		end
	end else begin
		for (i = 0; i < 16; i = i + 1) begin
			proposal_cnt[i] <= n_proposal_cnt[i];
		end
	end
end

always@* begin
    n_vid = vid_reg[batch_num_reg[3:0]]; // 16-1 mux
end

// dist_reg (checked)
always@(posedge clk) begin
    if(~rst_n_in) begin
        dist_reg <= 256'd0;
    end else begin
        dist_reg <= dist_rdata;
    end
end

// loc_oh_reg
always@(posedge clk) begin
    if(~rst_n_in) begin
        {loc_oh_reg[0], loc_oh_reg[1], loc_oh_reg[2], loc_oh_reg[3], loc_oh_reg[4], loc_oh_reg[5], loc_oh_reg[6], loc_oh_reg[7]} <= 128'd0;
        {loc_oh_reg[8], loc_oh_reg[9], loc_oh_reg[10], loc_oh_reg[11], loc_oh_reg[12], loc_oh_reg[13], loc_oh_reg[14], loc_oh_reg[15]} <= 128'd0;
        {loc_oh_reg[16], loc_oh_reg[17], loc_oh_reg[18], loc_oh_reg[19], loc_oh_reg[20], loc_oh_reg[21], loc_oh_reg[22], loc_oh_reg[23]} <= 128'd0;
        {loc_oh_reg[24], loc_oh_reg[25], loc_oh_reg[26], loc_oh_reg[27], loc_oh_reg[28], loc_oh_reg[29], loc_oh_reg[30], loc_oh_reg[31]} <= 128'd0;
        {loc_oh_reg[32], loc_oh_reg[33], loc_oh_reg[34], loc_oh_reg[35], loc_oh_reg[36], loc_oh_reg[37], loc_oh_reg[38], loc_oh_reg[39]} <= 128'd0;
        {loc_oh_reg[40], loc_oh_reg[41], loc_oh_reg[42], loc_oh_reg[43], loc_oh_reg[44], loc_oh_reg[45], loc_oh_reg[46], loc_oh_reg[47]} <= 128'd0;
        {loc_oh_reg[48], loc_oh_reg[49], loc_oh_reg[50], loc_oh_reg[51], loc_oh_reg[52], loc_oh_reg[53], loc_oh_reg[54], loc_oh_reg[55]} <= 128'd0;
        {loc_oh_reg[56], loc_oh_reg[57], loc_oh_reg[58], loc_oh_reg[59], loc_oh_reg[60], loc_oh_reg[61], loc_oh_reg[62], loc_oh_reg[63]} <= 128'd0;
        {loc_oh_reg[64], loc_oh_reg[65], loc_oh_reg[66], loc_oh_reg[67], loc_oh_reg[68], loc_oh_reg[69], loc_oh_reg[70], loc_oh_reg[71]} <= 128'd0;
        {loc_oh_reg[72], loc_oh_reg[73], loc_oh_reg[74], loc_oh_reg[75], loc_oh_reg[76], loc_oh_reg[77], loc_oh_reg[78], loc_oh_reg[79]} <= 128'd0;
        {loc_oh_reg[80], loc_oh_reg[81], loc_oh_reg[82], loc_oh_reg[83], loc_oh_reg[84], loc_oh_reg[85], loc_oh_reg[86], loc_oh_reg[87]} <= 128'd0;
        {loc_oh_reg[88], loc_oh_reg[89], loc_oh_reg[90], loc_oh_reg[91], loc_oh_reg[92], loc_oh_reg[93], loc_oh_reg[94], loc_oh_reg[95]} <= 128'd0;
        {loc_oh_reg[96], loc_oh_reg[97], loc_oh_reg[98], loc_oh_reg[99], loc_oh_reg[100], loc_oh_reg[101], loc_oh_reg[102], loc_oh_reg[103]} <= 128'd0;
        {loc_oh_reg[104], loc_oh_reg[105], loc_oh_reg[106], loc_oh_reg[107], loc_oh_reg[108], loc_oh_reg[109], loc_oh_reg[110], loc_oh_reg[111]} <= 128'd0;
        {loc_oh_reg[112], loc_oh_reg[113], loc_oh_reg[114], loc_oh_reg[115], loc_oh_reg[116], loc_oh_reg[117], loc_oh_reg[118], loc_oh_reg[119]} <= 128'd0;
        {loc_oh_reg[120], loc_oh_reg[121], loc_oh_reg[122], loc_oh_reg[123], loc_oh_reg[124], loc_oh_reg[125], loc_oh_reg[126], loc_oh_reg[127]} <= 128'd0;
        {loc_oh_reg[128], loc_oh_reg[129], loc_oh_reg[130], loc_oh_reg[131], loc_oh_reg[132], loc_oh_reg[133], loc_oh_reg[134], loc_oh_reg[135]} <= 128'd0;
        {loc_oh_reg[136], loc_oh_reg[137], loc_oh_reg[138], loc_oh_reg[139], loc_oh_reg[140], loc_oh_reg[141], loc_oh_reg[142], loc_oh_reg[143]} <= 128'd0;
        {loc_oh_reg[144], loc_oh_reg[145], loc_oh_reg[146], loc_oh_reg[147], loc_oh_reg[148], loc_oh_reg[149], loc_oh_reg[150], loc_oh_reg[151]} <= 128'd0;
        {loc_oh_reg[152], loc_oh_reg[153], loc_oh_reg[154], loc_oh_reg[155], loc_oh_reg[156], loc_oh_reg[157], loc_oh_reg[158], loc_oh_reg[159]} <= 128'd0;
        {loc_oh_reg[160], loc_oh_reg[161], loc_oh_reg[162], loc_oh_reg[163], loc_oh_reg[164], loc_oh_reg[165], loc_oh_reg[166], loc_oh_reg[167]} <= 128'd0;
        {loc_oh_reg[168], loc_oh_reg[169], loc_oh_reg[170], loc_oh_reg[171], loc_oh_reg[172], loc_oh_reg[173], loc_oh_reg[174], loc_oh_reg[175]} <= 128'd0;
        {loc_oh_reg[176], loc_oh_reg[177], loc_oh_reg[178], loc_oh_reg[179], loc_oh_reg[180], loc_oh_reg[181], loc_oh_reg[182], loc_oh_reg[183]} <= 128'd0;
        {loc_oh_reg[184], loc_oh_reg[185], loc_oh_reg[186], loc_oh_reg[187], loc_oh_reg[188], loc_oh_reg[189], loc_oh_reg[190], loc_oh_reg[191]} <= 128'd0;
        {loc_oh_reg[192], loc_oh_reg[193], loc_oh_reg[194], loc_oh_reg[195], loc_oh_reg[196], loc_oh_reg[197], loc_oh_reg[198], loc_oh_reg[199]} <= 128'd0;
        {loc_oh_reg[200], loc_oh_reg[201], loc_oh_reg[202], loc_oh_reg[203], loc_oh_reg[204], loc_oh_reg[205], loc_oh_reg[206], loc_oh_reg[207]} <= 128'd0;
        {loc_oh_reg[208], loc_oh_reg[209], loc_oh_reg[210], loc_oh_reg[211], loc_oh_reg[212], loc_oh_reg[213], loc_oh_reg[214], loc_oh_reg[215]} <= 128'd0;
        {loc_oh_reg[216], loc_oh_reg[217], loc_oh_reg[218], loc_oh_reg[219], loc_oh_reg[220], loc_oh_reg[221], loc_oh_reg[222], loc_oh_reg[223]} <= 128'd0;
        {loc_oh_reg[224], loc_oh_reg[225], loc_oh_reg[226], loc_oh_reg[227], loc_oh_reg[228], loc_oh_reg[229], loc_oh_reg[230], loc_oh_reg[231]} <= 128'd0;
        {loc_oh_reg[232], loc_oh_reg[233], loc_oh_reg[234], loc_oh_reg[235], loc_oh_reg[236], loc_oh_reg[237], loc_oh_reg[238], loc_oh_reg[239]} <= 128'd0;
        {loc_oh_reg[240], loc_oh_reg[241], loc_oh_reg[242], loc_oh_reg[243], loc_oh_reg[244], loc_oh_reg[245], loc_oh_reg[246], loc_oh_reg[247]} <= 128'd0;
        {loc_oh_reg[248], loc_oh_reg[249], loc_oh_reg[250], loc_oh_reg[251], loc_oh_reg[252], loc_oh_reg[253], loc_oh_reg[254], loc_oh_reg[255]} <= 128'd0;
    end else begin
        {loc_oh_reg[0], loc_oh_reg[1], loc_oh_reg[2], loc_oh_reg[3], loc_oh_reg[4], loc_oh_reg[5], loc_oh_reg[6], loc_oh_reg[7]} <= {n_loc_oh_reg[0], n_loc_oh_reg[1], n_loc_oh_reg[2], n_loc_oh_reg[3], n_loc_oh_reg[4], n_loc_oh_reg[5], n_loc_oh_reg[6], n_loc_oh_reg[7]};
        {loc_oh_reg[8], loc_oh_reg[9], loc_oh_reg[10], loc_oh_reg[11], loc_oh_reg[12], loc_oh_reg[13], loc_oh_reg[14], loc_oh_reg[15]} <= {n_loc_oh_reg[8], n_loc_oh_reg[9], n_loc_oh_reg[10], n_loc_oh_reg[11], n_loc_oh_reg[12], n_loc_oh_reg[13], n_loc_oh_reg[14], n_loc_oh_reg[15]};
        {loc_oh_reg[16], loc_oh_reg[17], loc_oh_reg[18], loc_oh_reg[19], loc_oh_reg[20], loc_oh_reg[21], loc_oh_reg[22], loc_oh_reg[23]} <= {n_loc_oh_reg[16], n_loc_oh_reg[17], n_loc_oh_reg[18], n_loc_oh_reg[19], n_loc_oh_reg[20], n_loc_oh_reg[21], n_loc_oh_reg[22], n_loc_oh_reg[23]};
        {loc_oh_reg[24], loc_oh_reg[25], loc_oh_reg[26], loc_oh_reg[27], loc_oh_reg[28], loc_oh_reg[29], loc_oh_reg[30], loc_oh_reg[31]} <= {n_loc_oh_reg[24], n_loc_oh_reg[25], n_loc_oh_reg[26], n_loc_oh_reg[27], n_loc_oh_reg[28], n_loc_oh_reg[29], n_loc_oh_reg[30], n_loc_oh_reg[31]};
        {loc_oh_reg[32], loc_oh_reg[33], loc_oh_reg[34], loc_oh_reg[35], loc_oh_reg[36], loc_oh_reg[37], loc_oh_reg[38], loc_oh_reg[39]} <= {n_loc_oh_reg[32], n_loc_oh_reg[33], n_loc_oh_reg[34], n_loc_oh_reg[35], n_loc_oh_reg[36], n_loc_oh_reg[37], n_loc_oh_reg[38], n_loc_oh_reg[39]};
        {loc_oh_reg[40], loc_oh_reg[41], loc_oh_reg[42], loc_oh_reg[43], loc_oh_reg[44], loc_oh_reg[45], loc_oh_reg[46], loc_oh_reg[47]} <= {n_loc_oh_reg[40], n_loc_oh_reg[41], n_loc_oh_reg[42], n_loc_oh_reg[43], n_loc_oh_reg[44], n_loc_oh_reg[45], n_loc_oh_reg[46], n_loc_oh_reg[47]};
        {loc_oh_reg[48], loc_oh_reg[49], loc_oh_reg[50], loc_oh_reg[51], loc_oh_reg[52], loc_oh_reg[53], loc_oh_reg[54], loc_oh_reg[55]} <= {n_loc_oh_reg[48], n_loc_oh_reg[49], n_loc_oh_reg[50], n_loc_oh_reg[51], n_loc_oh_reg[52], n_loc_oh_reg[53], n_loc_oh_reg[54], n_loc_oh_reg[55]};
        {loc_oh_reg[56], loc_oh_reg[57], loc_oh_reg[58], loc_oh_reg[59], loc_oh_reg[60], loc_oh_reg[61], loc_oh_reg[62], loc_oh_reg[63]} <= {n_loc_oh_reg[56], n_loc_oh_reg[57], n_loc_oh_reg[58], n_loc_oh_reg[59], n_loc_oh_reg[60], n_loc_oh_reg[61], n_loc_oh_reg[62], n_loc_oh_reg[63]};
        {loc_oh_reg[64], loc_oh_reg[65], loc_oh_reg[66], loc_oh_reg[67], loc_oh_reg[68], loc_oh_reg[69], loc_oh_reg[70], loc_oh_reg[71]} <= {n_loc_oh_reg[64], n_loc_oh_reg[65], n_loc_oh_reg[66], n_loc_oh_reg[67], n_loc_oh_reg[68], n_loc_oh_reg[69], n_loc_oh_reg[70], n_loc_oh_reg[71]};
        {loc_oh_reg[72], loc_oh_reg[73], loc_oh_reg[74], loc_oh_reg[75], loc_oh_reg[76], loc_oh_reg[77], loc_oh_reg[78], loc_oh_reg[79]} <= {n_loc_oh_reg[72], n_loc_oh_reg[73], n_loc_oh_reg[74], n_loc_oh_reg[75], n_loc_oh_reg[76], n_loc_oh_reg[77], n_loc_oh_reg[78], n_loc_oh_reg[79]};
        {loc_oh_reg[80], loc_oh_reg[81], loc_oh_reg[82], loc_oh_reg[83], loc_oh_reg[84], loc_oh_reg[85], loc_oh_reg[86], loc_oh_reg[87]} <= {n_loc_oh_reg[80], n_loc_oh_reg[81], n_loc_oh_reg[82], n_loc_oh_reg[83], n_loc_oh_reg[84], n_loc_oh_reg[85], n_loc_oh_reg[86], n_loc_oh_reg[87]};
        {loc_oh_reg[88], loc_oh_reg[89], loc_oh_reg[90], loc_oh_reg[91], loc_oh_reg[92], loc_oh_reg[93], loc_oh_reg[94], loc_oh_reg[95]} <= {n_loc_oh_reg[88], n_loc_oh_reg[89], n_loc_oh_reg[90], n_loc_oh_reg[91], n_loc_oh_reg[92], n_loc_oh_reg[93], n_loc_oh_reg[94], n_loc_oh_reg[95]};
        {loc_oh_reg[96], loc_oh_reg[97], loc_oh_reg[98], loc_oh_reg[99], loc_oh_reg[100], loc_oh_reg[101], loc_oh_reg[102], loc_oh_reg[103]} <= {n_loc_oh_reg[96], n_loc_oh_reg[97], n_loc_oh_reg[98], n_loc_oh_reg[99], n_loc_oh_reg[100], n_loc_oh_reg[101], n_loc_oh_reg[102], n_loc_oh_reg[103]};
        {loc_oh_reg[104], loc_oh_reg[105], loc_oh_reg[106], loc_oh_reg[107], loc_oh_reg[108], loc_oh_reg[109], loc_oh_reg[110], loc_oh_reg[111]} <= {n_loc_oh_reg[104], n_loc_oh_reg[105], n_loc_oh_reg[106], n_loc_oh_reg[107], n_loc_oh_reg[108], n_loc_oh_reg[109], n_loc_oh_reg[110], n_loc_oh_reg[111]};
        {loc_oh_reg[112], loc_oh_reg[113], loc_oh_reg[114], loc_oh_reg[115], loc_oh_reg[116], loc_oh_reg[117], loc_oh_reg[118], loc_oh_reg[119]} <= {n_loc_oh_reg[112], n_loc_oh_reg[113], n_loc_oh_reg[114], n_loc_oh_reg[115], n_loc_oh_reg[116], n_loc_oh_reg[117], n_loc_oh_reg[118], n_loc_oh_reg[119]};
        {loc_oh_reg[120], loc_oh_reg[121], loc_oh_reg[122], loc_oh_reg[123], loc_oh_reg[124], loc_oh_reg[125], loc_oh_reg[126], loc_oh_reg[127]} <= {n_loc_oh_reg[120], n_loc_oh_reg[121], n_loc_oh_reg[122], n_loc_oh_reg[123], n_loc_oh_reg[124], n_loc_oh_reg[125], n_loc_oh_reg[126], n_loc_oh_reg[127]};
        {loc_oh_reg[128], loc_oh_reg[129], loc_oh_reg[130], loc_oh_reg[131], loc_oh_reg[132], loc_oh_reg[133], loc_oh_reg[134], loc_oh_reg[135]} <= {n_loc_oh_reg[128], n_loc_oh_reg[129], n_loc_oh_reg[130], n_loc_oh_reg[131], n_loc_oh_reg[132], n_loc_oh_reg[133], n_loc_oh_reg[134], n_loc_oh_reg[135]};
        {loc_oh_reg[136], loc_oh_reg[137], loc_oh_reg[138], loc_oh_reg[139], loc_oh_reg[140], loc_oh_reg[141], loc_oh_reg[142], loc_oh_reg[143]} <= {n_loc_oh_reg[136], n_loc_oh_reg[137], n_loc_oh_reg[138], n_loc_oh_reg[139], n_loc_oh_reg[140], n_loc_oh_reg[141], n_loc_oh_reg[142], n_loc_oh_reg[143]};
        {loc_oh_reg[144], loc_oh_reg[145], loc_oh_reg[146], loc_oh_reg[147], loc_oh_reg[148], loc_oh_reg[149], loc_oh_reg[150], loc_oh_reg[151]} <= {n_loc_oh_reg[144], n_loc_oh_reg[145], n_loc_oh_reg[146], n_loc_oh_reg[147], n_loc_oh_reg[148], n_loc_oh_reg[149], n_loc_oh_reg[150], n_loc_oh_reg[151]};
        {loc_oh_reg[152], loc_oh_reg[153], loc_oh_reg[154], loc_oh_reg[155], loc_oh_reg[156], loc_oh_reg[157], loc_oh_reg[158], loc_oh_reg[159]} <= {n_loc_oh_reg[152], n_loc_oh_reg[153], n_loc_oh_reg[154], n_loc_oh_reg[155], n_loc_oh_reg[156], n_loc_oh_reg[157], n_loc_oh_reg[158], n_loc_oh_reg[159]};
        {loc_oh_reg[160], loc_oh_reg[161], loc_oh_reg[162], loc_oh_reg[163], loc_oh_reg[164], loc_oh_reg[165], loc_oh_reg[166], loc_oh_reg[167]} <= {n_loc_oh_reg[160], n_loc_oh_reg[161], n_loc_oh_reg[162], n_loc_oh_reg[163], n_loc_oh_reg[164], n_loc_oh_reg[165], n_loc_oh_reg[166], n_loc_oh_reg[167]};
        {loc_oh_reg[168], loc_oh_reg[169], loc_oh_reg[170], loc_oh_reg[171], loc_oh_reg[172], loc_oh_reg[173], loc_oh_reg[174], loc_oh_reg[175]} <= {n_loc_oh_reg[168], n_loc_oh_reg[169], n_loc_oh_reg[170], n_loc_oh_reg[171], n_loc_oh_reg[172], n_loc_oh_reg[173], n_loc_oh_reg[174], n_loc_oh_reg[175]};
        {loc_oh_reg[176], loc_oh_reg[177], loc_oh_reg[178], loc_oh_reg[179], loc_oh_reg[180], loc_oh_reg[181], loc_oh_reg[182], loc_oh_reg[183]} <= {n_loc_oh_reg[176], n_loc_oh_reg[177], n_loc_oh_reg[178], n_loc_oh_reg[179], n_loc_oh_reg[180], n_loc_oh_reg[181], n_loc_oh_reg[182], n_loc_oh_reg[183]};
        {loc_oh_reg[184], loc_oh_reg[185], loc_oh_reg[186], loc_oh_reg[187], loc_oh_reg[188], loc_oh_reg[189], loc_oh_reg[190], loc_oh_reg[191]} <= {n_loc_oh_reg[184], n_loc_oh_reg[185], n_loc_oh_reg[186], n_loc_oh_reg[187], n_loc_oh_reg[188], n_loc_oh_reg[189], n_loc_oh_reg[190], n_loc_oh_reg[191]};
        {loc_oh_reg[192], loc_oh_reg[193], loc_oh_reg[194], loc_oh_reg[195], loc_oh_reg[196], loc_oh_reg[197], loc_oh_reg[198], loc_oh_reg[199]} <= {n_loc_oh_reg[192], n_loc_oh_reg[193], n_loc_oh_reg[194], n_loc_oh_reg[195], n_loc_oh_reg[196], n_loc_oh_reg[197], n_loc_oh_reg[198], n_loc_oh_reg[199]};
        {loc_oh_reg[200], loc_oh_reg[201], loc_oh_reg[202], loc_oh_reg[203], loc_oh_reg[204], loc_oh_reg[205], loc_oh_reg[206], loc_oh_reg[207]} <= {n_loc_oh_reg[200], n_loc_oh_reg[201], n_loc_oh_reg[202], n_loc_oh_reg[203], n_loc_oh_reg[204], n_loc_oh_reg[205], n_loc_oh_reg[206], n_loc_oh_reg[207]};
        {loc_oh_reg[208], loc_oh_reg[209], loc_oh_reg[210], loc_oh_reg[211], loc_oh_reg[212], loc_oh_reg[213], loc_oh_reg[214], loc_oh_reg[215]} <= {n_loc_oh_reg[208], n_loc_oh_reg[209], n_loc_oh_reg[210], n_loc_oh_reg[211], n_loc_oh_reg[212], n_loc_oh_reg[213], n_loc_oh_reg[214], n_loc_oh_reg[215]};
        {loc_oh_reg[216], loc_oh_reg[217], loc_oh_reg[218], loc_oh_reg[219], loc_oh_reg[220], loc_oh_reg[221], loc_oh_reg[222], loc_oh_reg[223]} <= {n_loc_oh_reg[216], n_loc_oh_reg[217], n_loc_oh_reg[218], n_loc_oh_reg[219], n_loc_oh_reg[220], n_loc_oh_reg[221], n_loc_oh_reg[222], n_loc_oh_reg[223]};
        {loc_oh_reg[224], loc_oh_reg[225], loc_oh_reg[226], loc_oh_reg[227], loc_oh_reg[228], loc_oh_reg[229], loc_oh_reg[230], loc_oh_reg[231]} <= {n_loc_oh_reg[224], n_loc_oh_reg[225], n_loc_oh_reg[226], n_loc_oh_reg[227], n_loc_oh_reg[228], n_loc_oh_reg[229], n_loc_oh_reg[230], n_loc_oh_reg[231]};
        {loc_oh_reg[232], loc_oh_reg[233], loc_oh_reg[234], loc_oh_reg[235], loc_oh_reg[236], loc_oh_reg[237], loc_oh_reg[238], loc_oh_reg[239]} <= {n_loc_oh_reg[232], n_loc_oh_reg[233], n_loc_oh_reg[234], n_loc_oh_reg[235], n_loc_oh_reg[236], n_loc_oh_reg[237], n_loc_oh_reg[238], n_loc_oh_reg[239]};
        {loc_oh_reg[240], loc_oh_reg[241], loc_oh_reg[242], loc_oh_reg[243], loc_oh_reg[244], loc_oh_reg[245], loc_oh_reg[246], loc_oh_reg[247]} <= {n_loc_oh_reg[240], n_loc_oh_reg[241], n_loc_oh_reg[242], n_loc_oh_reg[243], n_loc_oh_reg[244], n_loc_oh_reg[245], n_loc_oh_reg[246], n_loc_oh_reg[247]};
        {loc_oh_reg[248], loc_oh_reg[249], loc_oh_reg[250], loc_oh_reg[251], loc_oh_reg[252], loc_oh_reg[253], loc_oh_reg[254], loc_oh_reg[255]} <= {n_loc_oh_reg[248], n_loc_oh_reg[249], n_loc_oh_reg[250], n_loc_oh_reg[251], n_loc_oh_reg[252], n_loc_oh_reg[253], n_loc_oh_reg[254], n_loc_oh_reg[255]};
    end
end

// dsum
always@(posedge clk) begin
    if(~rst_n_in) begin
        {dsum_reg[0], dsum_reg[1], dsum_reg[2], dsum_reg[3], dsum_reg[4], dsum_reg[5], dsum_reg[6], dsum_reg[7]} <= 40'd0;
        {dsum_reg[8], dsum_reg[9], dsum_reg[10], dsum_reg[11], dsum_reg[12], dsum_reg[13], dsum_reg[14], dsum_reg[15]} <= 40'd0;
        {dsum_reg[16], dsum_reg[17], dsum_reg[18], dsum_reg[19], dsum_reg[20], dsum_reg[21], dsum_reg[22], dsum_reg[23]} <= 40'd0;
        {dsum_reg[24], dsum_reg[25], dsum_reg[26], dsum_reg[27], dsum_reg[28], dsum_reg[29], dsum_reg[30], dsum_reg[31]} <= 40'd0;
        {dsum_reg[32], dsum_reg[33], dsum_reg[34], dsum_reg[35], dsum_reg[36], dsum_reg[37], dsum_reg[38], dsum_reg[39]} <= 40'd0;
        {dsum_reg[40], dsum_reg[41], dsum_reg[42], dsum_reg[43], dsum_reg[44], dsum_reg[45], dsum_reg[46], dsum_reg[47]} <= 40'd0;
        {dsum_reg[48], dsum_reg[49], dsum_reg[50], dsum_reg[51], dsum_reg[52], dsum_reg[53], dsum_reg[54], dsum_reg[55]} <= 40'd0;
        {dsum_reg[56], dsum_reg[57], dsum_reg[58], dsum_reg[59], dsum_reg[60], dsum_reg[61], dsum_reg[62], dsum_reg[63]} <= 40'd0;
        {dsum_reg[64], dsum_reg[65], dsum_reg[66], dsum_reg[67], dsum_reg[68], dsum_reg[69], dsum_reg[70], dsum_reg[71]} <= 40'd0;
        {dsum_reg[72], dsum_reg[73], dsum_reg[74], dsum_reg[75], dsum_reg[76], dsum_reg[77], dsum_reg[78], dsum_reg[79]} <= 40'd0;
        {dsum_reg[80], dsum_reg[81], dsum_reg[82], dsum_reg[83], dsum_reg[84], dsum_reg[85], dsum_reg[86], dsum_reg[87]} <= 40'd0;
        {dsum_reg[88], dsum_reg[89], dsum_reg[90], dsum_reg[91], dsum_reg[92], dsum_reg[93], dsum_reg[94], dsum_reg[95]} <= 40'd0;
        {dsum_reg[96], dsum_reg[97], dsum_reg[98], dsum_reg[99], dsum_reg[100], dsum_reg[101], dsum_reg[102], dsum_reg[103]} <= 40'd0;
        {dsum_reg[104], dsum_reg[105], dsum_reg[106], dsum_reg[107], dsum_reg[108], dsum_reg[109], dsum_reg[110], dsum_reg[111]} <= 40'd0;
        {dsum_reg[112], dsum_reg[113], dsum_reg[114], dsum_reg[115], dsum_reg[116], dsum_reg[117], dsum_reg[118], dsum_reg[119]} <= 40'd0;
        {dsum_reg[120], dsum_reg[121], dsum_reg[122], dsum_reg[123], dsum_reg[124], dsum_reg[125], dsum_reg[126], dsum_reg[127]} <= 40'd0;
    end else begin
        {dsum_reg[0], dsum_reg[1], dsum_reg[2], dsum_reg[3], dsum_reg[4], dsum_reg[5], dsum_reg[6], dsum_reg[7]} <= {n_dsum_reg[0], n_dsum_reg[1], n_dsum_reg[2], n_dsum_reg[3], n_dsum_reg[4], n_dsum_reg[5], n_dsum_reg[6], n_dsum_reg[7]};
        {dsum_reg[8], dsum_reg[9], dsum_reg[10], dsum_reg[11], dsum_reg[12], dsum_reg[13], dsum_reg[14], dsum_reg[15]} <= {n_dsum_reg[8], n_dsum_reg[9], n_dsum_reg[10], n_dsum_reg[11], n_dsum_reg[12], n_dsum_reg[13], n_dsum_reg[14], n_dsum_reg[15]};
        {dsum_reg[16], dsum_reg[17], dsum_reg[18], dsum_reg[19], dsum_reg[20], dsum_reg[21], dsum_reg[22], dsum_reg[23]} <= {n_dsum_reg[16], n_dsum_reg[17], n_dsum_reg[18], n_dsum_reg[19], n_dsum_reg[20], n_dsum_reg[21], n_dsum_reg[22], n_dsum_reg[23]};
        {dsum_reg[24], dsum_reg[25], dsum_reg[26], dsum_reg[27], dsum_reg[28], dsum_reg[29], dsum_reg[30], dsum_reg[31]} <= {n_dsum_reg[24], n_dsum_reg[25], n_dsum_reg[26], n_dsum_reg[27], n_dsum_reg[28], n_dsum_reg[29], n_dsum_reg[30], n_dsum_reg[31]};
        {dsum_reg[32], dsum_reg[33], dsum_reg[34], dsum_reg[35], dsum_reg[36], dsum_reg[37], dsum_reg[38], dsum_reg[39]} <= {n_dsum_reg[32], n_dsum_reg[33], n_dsum_reg[34], n_dsum_reg[35], n_dsum_reg[36], n_dsum_reg[37], n_dsum_reg[38], n_dsum_reg[39]};
        {dsum_reg[40], dsum_reg[41], dsum_reg[42], dsum_reg[43], dsum_reg[44], dsum_reg[45], dsum_reg[46], dsum_reg[47]} <= {n_dsum_reg[40], n_dsum_reg[41], n_dsum_reg[42], n_dsum_reg[43], n_dsum_reg[44], n_dsum_reg[45], n_dsum_reg[46], n_dsum_reg[47]};
        {dsum_reg[48], dsum_reg[49], dsum_reg[50], dsum_reg[51], dsum_reg[52], dsum_reg[53], dsum_reg[54], dsum_reg[55]} <= {n_dsum_reg[48], n_dsum_reg[49], n_dsum_reg[50], n_dsum_reg[51], n_dsum_reg[52], n_dsum_reg[53], n_dsum_reg[54], n_dsum_reg[55]};
        {dsum_reg[56], dsum_reg[57], dsum_reg[58], dsum_reg[59], dsum_reg[60], dsum_reg[61], dsum_reg[62], dsum_reg[63]} <= {n_dsum_reg[56], n_dsum_reg[57], n_dsum_reg[58], n_dsum_reg[59], n_dsum_reg[60], n_dsum_reg[61], n_dsum_reg[62], n_dsum_reg[63]};
        {dsum_reg[64], dsum_reg[65], dsum_reg[66], dsum_reg[67], dsum_reg[68], dsum_reg[69], dsum_reg[70], dsum_reg[71]} <= {n_dsum_reg[64], n_dsum_reg[65], n_dsum_reg[66], n_dsum_reg[67], n_dsum_reg[68], n_dsum_reg[69], n_dsum_reg[70], n_dsum_reg[71]};
        {dsum_reg[72], dsum_reg[73], dsum_reg[74], dsum_reg[75], dsum_reg[76], dsum_reg[77], dsum_reg[78], dsum_reg[79]} <= {n_dsum_reg[72], n_dsum_reg[73], n_dsum_reg[74], n_dsum_reg[75], n_dsum_reg[76], n_dsum_reg[77], n_dsum_reg[78], n_dsum_reg[79]};
        {dsum_reg[80], dsum_reg[81], dsum_reg[82], dsum_reg[83], dsum_reg[84], dsum_reg[85], dsum_reg[86], dsum_reg[87]} <= {n_dsum_reg[80], n_dsum_reg[81], n_dsum_reg[82], n_dsum_reg[83], n_dsum_reg[84], n_dsum_reg[85], n_dsum_reg[86], n_dsum_reg[87]};
        {dsum_reg[88], dsum_reg[89], dsum_reg[90], dsum_reg[91], dsum_reg[92], dsum_reg[93], dsum_reg[94], dsum_reg[95]} <= {n_dsum_reg[88], n_dsum_reg[89], n_dsum_reg[90], n_dsum_reg[91], n_dsum_reg[92], n_dsum_reg[93], n_dsum_reg[94], n_dsum_reg[95]};
        {dsum_reg[96], dsum_reg[97], dsum_reg[98], dsum_reg[99], dsum_reg[100], dsum_reg[101], dsum_reg[102], dsum_reg[103]} <= {n_dsum_reg[96], n_dsum_reg[97], n_dsum_reg[98], n_dsum_reg[99], n_dsum_reg[100], n_dsum_reg[101], n_dsum_reg[102], n_dsum_reg[103]};
        {dsum_reg[104], dsum_reg[105], dsum_reg[106], dsum_reg[107], dsum_reg[108], dsum_reg[109], dsum_reg[110], dsum_reg[111]} <= {n_dsum_reg[104], n_dsum_reg[105], n_dsum_reg[106], n_dsum_reg[107], n_dsum_reg[108], n_dsum_reg[109], n_dsum_reg[110], n_dsum_reg[111]};
        {dsum_reg[112], dsum_reg[113], dsum_reg[114], dsum_reg[115], dsum_reg[116], dsum_reg[117], dsum_reg[118], dsum_reg[119]} <= {n_dsum_reg[112], n_dsum_reg[113], n_dsum_reg[114], n_dsum_reg[115], n_dsum_reg[116], n_dsum_reg[117], n_dsum_reg[118], n_dsum_reg[119]};
        {dsum_reg[120], dsum_reg[121], dsum_reg[122], dsum_reg[123], dsum_reg[124], dsum_reg[125], dsum_reg[126], dsum_reg[127]} <= {n_dsum_reg[120], n_dsum_reg[121], n_dsum_reg[122], n_dsum_reg[123], n_dsum_reg[124], n_dsum_reg[125], n_dsum_reg[126], n_dsum_reg[127]};
    end
end

// part
always@(posedge clk) begin
    if(~rst_n_in) begin
        {part_reg[0], part_reg[1], part_reg[2], part_reg[3], part_reg[4], part_reg[5], part_reg[6], part_reg[7]} <= 32'd0;
        {part_reg[8], part_reg[9], part_reg[10], part_reg[11], part_reg[12], part_reg[13], part_reg[14], part_reg[15]} <= 32'd0;
    end else begin
        {part_reg[0], part_reg[1], part_reg[2], part_reg[3], part_reg[4], part_reg[5], part_reg[6], part_reg[7]} <= {n_part_reg[0], n_part_reg[1], n_part_reg[2], n_part_reg[3], n_part_reg[4], n_part_reg[5], n_part_reg[6], n_part_reg[7]};
        {part_reg[8], part_reg[9], part_reg[10], part_reg[11], part_reg[12], part_reg[13], part_reg[14], part_reg[15]} <= {n_part_reg[8], n_part_reg[9], n_part_reg[10], n_part_reg[11], n_part_reg[12], n_part_reg[13], n_part_reg[14], n_part_reg[15]};
    end
end

// loc_reg (checked)
always@(posedge clk) begin
    if(~rst_n_in) begin
        {loc_reg[0], loc_reg[1], loc_reg[2], loc_reg[3], loc_reg[4], loc_reg[5], loc_reg[6], loc_reg[7]} <= 32'd0;
        {loc_reg[8], loc_reg[9], loc_reg[10], loc_reg[11], loc_reg[12], loc_reg[13], loc_reg[14], loc_reg[15]} <= 32'd0;
        {loc_reg[16], loc_reg[17], loc_reg[18], loc_reg[19], loc_reg[20], loc_reg[21], loc_reg[22], loc_reg[23]} <= 32'd0;
        {loc_reg[24], loc_reg[25], loc_reg[26], loc_reg[27], loc_reg[28], loc_reg[29], loc_reg[30], loc_reg[31]} <= 32'd0;
        {loc_reg[32], loc_reg[33], loc_reg[34], loc_reg[35], loc_reg[36], loc_reg[37], loc_reg[38], loc_reg[39]} <= 32'd0;
        {loc_reg[40], loc_reg[41], loc_reg[42], loc_reg[43], loc_reg[44], loc_reg[45], loc_reg[46], loc_reg[47]} <= 32'd0;
        {loc_reg[48], loc_reg[49], loc_reg[50], loc_reg[51], loc_reg[52], loc_reg[53], loc_reg[54], loc_reg[55]} <= 32'd0;
        {loc_reg[56], loc_reg[57], loc_reg[58], loc_reg[59], loc_reg[60], loc_reg[61], loc_reg[62], loc_reg[63]} <= 32'd0;
        {loc_reg[64], loc_reg[65], loc_reg[66], loc_reg[67], loc_reg[68], loc_reg[69], loc_reg[70], loc_reg[71]} <= 32'd0;
        {loc_reg[72], loc_reg[73], loc_reg[74], loc_reg[75], loc_reg[76], loc_reg[77], loc_reg[78], loc_reg[79]} <= 32'd0;
        {loc_reg[80], loc_reg[81], loc_reg[82], loc_reg[83], loc_reg[84], loc_reg[85], loc_reg[86], loc_reg[87]} <= 32'd0;
        {loc_reg[88], loc_reg[89], loc_reg[90], loc_reg[91], loc_reg[92], loc_reg[93], loc_reg[94], loc_reg[95]} <= 32'd0;
        {loc_reg[96], loc_reg[97], loc_reg[98], loc_reg[99], loc_reg[100], loc_reg[101], loc_reg[102], loc_reg[103]} <= 32'd0;
        {loc_reg[104], loc_reg[105], loc_reg[106], loc_reg[107], loc_reg[108], loc_reg[109], loc_reg[110], loc_reg[111]} <= 32'd0;
        {loc_reg[112], loc_reg[113], loc_reg[114], loc_reg[115], loc_reg[116], loc_reg[117], loc_reg[118], loc_reg[119]} <= 32'd0;
        {loc_reg[120], loc_reg[121], loc_reg[122], loc_reg[123], loc_reg[124], loc_reg[125], loc_reg[126], loc_reg[127]} <= 32'd0;
        {loc_reg[128], loc_reg[129], loc_reg[130], loc_reg[131], loc_reg[132], loc_reg[133], loc_reg[134], loc_reg[135]} <= 32'd0;
        {loc_reg[136], loc_reg[137], loc_reg[138], loc_reg[139], loc_reg[140], loc_reg[141], loc_reg[142], loc_reg[143]} <= 32'd0;
        {loc_reg[144], loc_reg[145], loc_reg[146], loc_reg[147], loc_reg[148], loc_reg[149], loc_reg[150], loc_reg[151]} <= 32'd0;
        {loc_reg[152], loc_reg[153], loc_reg[154], loc_reg[155], loc_reg[156], loc_reg[157], loc_reg[158], loc_reg[159]} <= 32'd0;
        {loc_reg[160], loc_reg[161], loc_reg[162], loc_reg[163], loc_reg[164], loc_reg[165], loc_reg[166], loc_reg[167]} <= 32'd0;
        {loc_reg[168], loc_reg[169], loc_reg[170], loc_reg[171], loc_reg[172], loc_reg[173], loc_reg[174], loc_reg[175]} <= 32'd0;
        {loc_reg[176], loc_reg[177], loc_reg[178], loc_reg[179], loc_reg[180], loc_reg[181], loc_reg[182], loc_reg[183]} <= 32'd0;
        {loc_reg[184], loc_reg[185], loc_reg[186], loc_reg[187], loc_reg[188], loc_reg[189], loc_reg[190], loc_reg[191]} <= 32'd0;
        {loc_reg[192], loc_reg[193], loc_reg[194], loc_reg[195], loc_reg[196], loc_reg[197], loc_reg[198], loc_reg[199]} <= 32'd0;
        {loc_reg[200], loc_reg[201], loc_reg[202], loc_reg[203], loc_reg[204], loc_reg[205], loc_reg[206], loc_reg[207]} <= 32'd0;
        {loc_reg[208], loc_reg[209], loc_reg[210], loc_reg[211], loc_reg[212], loc_reg[213], loc_reg[214], loc_reg[215]} <= 32'd0;
        {loc_reg[216], loc_reg[217], loc_reg[218], loc_reg[219], loc_reg[220], loc_reg[221], loc_reg[222], loc_reg[223]} <= 32'd0;
        {loc_reg[224], loc_reg[225], loc_reg[226], loc_reg[227], loc_reg[228], loc_reg[229], loc_reg[230], loc_reg[231]} <= 32'd0;
        {loc_reg[232], loc_reg[233], loc_reg[234], loc_reg[235], loc_reg[236], loc_reg[237], loc_reg[238], loc_reg[239]} <= 32'd0;
        {loc_reg[240], loc_reg[241], loc_reg[242], loc_reg[243], loc_reg[244], loc_reg[245], loc_reg[246], loc_reg[247]} <= 32'd0;
        {loc_reg[248], loc_reg[249], loc_reg[250], loc_reg[251], loc_reg[252], loc_reg[253], loc_reg[254], loc_reg[255]} <= 32'd0;
    end else begin
        {loc_reg[0], loc_reg[1], loc_reg[2], loc_reg[3], loc_reg[4], loc_reg[5], loc_reg[6], loc_reg[7]} <= {loc_rdata[1023:1020], loc_rdata[1019:1016], loc_rdata[1015:1012], loc_rdata[1011:1008], loc_rdata[1007:1004], loc_rdata[1003:1000], loc_rdata[999:996], loc_rdata[995:992]};
        {loc_reg[8], loc_reg[9], loc_reg[10], loc_reg[11], loc_reg[12], loc_reg[13], loc_reg[14], loc_reg[15]} <= {loc_rdata[991:988], loc_rdata[987:984], loc_rdata[983:980], loc_rdata[979:976], loc_rdata[975:972], loc_rdata[971:968], loc_rdata[967:964], loc_rdata[963:960]};
        {loc_reg[16], loc_reg[17], loc_reg[18], loc_reg[19], loc_reg[20], loc_reg[21], loc_reg[22], loc_reg[23]} <= {loc_rdata[959:956], loc_rdata[955:952], loc_rdata[951:948], loc_rdata[947:944], loc_rdata[943:940], loc_rdata[939:936], loc_rdata[935:932], loc_rdata[931:928]};
        {loc_reg[24], loc_reg[25], loc_reg[26], loc_reg[27], loc_reg[28], loc_reg[29], loc_reg[30], loc_reg[31]} <= {loc_rdata[927:924], loc_rdata[923:920], loc_rdata[919:916], loc_rdata[915:912], loc_rdata[911:908], loc_rdata[907:904], loc_rdata[903:900], loc_rdata[899:896]};
        {loc_reg[32], loc_reg[33], loc_reg[34], loc_reg[35], loc_reg[36], loc_reg[37], loc_reg[38], loc_reg[39]} <= {loc_rdata[895:892], loc_rdata[891:888], loc_rdata[887:884], loc_rdata[883:880], loc_rdata[879:876], loc_rdata[875:872], loc_rdata[871:868], loc_rdata[867:864]};
        {loc_reg[40], loc_reg[41], loc_reg[42], loc_reg[43], loc_reg[44], loc_reg[45], loc_reg[46], loc_reg[47]} <= {loc_rdata[863:860], loc_rdata[859:856], loc_rdata[855:852], loc_rdata[851:848], loc_rdata[847:844], loc_rdata[843:840], loc_rdata[839:836], loc_rdata[835:832]};
        {loc_reg[48], loc_reg[49], loc_reg[50], loc_reg[51], loc_reg[52], loc_reg[53], loc_reg[54], loc_reg[55]} <= {loc_rdata[831:828], loc_rdata[827:824], loc_rdata[823:820], loc_rdata[819:816], loc_rdata[815:812], loc_rdata[811:808], loc_rdata[807:804], loc_rdata[803:800]};
        {loc_reg[56], loc_reg[57], loc_reg[58], loc_reg[59], loc_reg[60], loc_reg[61], loc_reg[62], loc_reg[63]} <= {loc_rdata[799:796], loc_rdata[795:792], loc_rdata[791:788], loc_rdata[787:784], loc_rdata[783:780], loc_rdata[779:776], loc_rdata[775:772], loc_rdata[771:768]};
        {loc_reg[64], loc_reg[65], loc_reg[66], loc_reg[67], loc_reg[68], loc_reg[69], loc_reg[70], loc_reg[71]} <= {loc_rdata[767:764], loc_rdata[763:760], loc_rdata[759:756], loc_rdata[755:752], loc_rdata[751:748], loc_rdata[747:744], loc_rdata[743:740], loc_rdata[739:736]};
        {loc_reg[72], loc_reg[73], loc_reg[74], loc_reg[75], loc_reg[76], loc_reg[77], loc_reg[78], loc_reg[79]} <= {loc_rdata[735:732], loc_rdata[731:728], loc_rdata[727:724], loc_rdata[723:720], loc_rdata[719:716], loc_rdata[715:712], loc_rdata[711:708], loc_rdata[707:704]};
        {loc_reg[80], loc_reg[81], loc_reg[82], loc_reg[83], loc_reg[84], loc_reg[85], loc_reg[86], loc_reg[87]} <= {loc_rdata[703:700], loc_rdata[699:696], loc_rdata[695:692], loc_rdata[691:688], loc_rdata[687:684], loc_rdata[683:680], loc_rdata[679:676], loc_rdata[675:672]};
        {loc_reg[88], loc_reg[89], loc_reg[90], loc_reg[91], loc_reg[92], loc_reg[93], loc_reg[94], loc_reg[95]} <= {loc_rdata[671:668], loc_rdata[667:664], loc_rdata[663:660], loc_rdata[659:656], loc_rdata[655:652], loc_rdata[651:648], loc_rdata[647:644], loc_rdata[643:640]};
        {loc_reg[96], loc_reg[97], loc_reg[98], loc_reg[99], loc_reg[100], loc_reg[101], loc_reg[102], loc_reg[103]} <= {loc_rdata[639:636], loc_rdata[635:632], loc_rdata[631:628], loc_rdata[627:624], loc_rdata[623:620], loc_rdata[619:616], loc_rdata[615:612], loc_rdata[611:608]};
        {loc_reg[104], loc_reg[105], loc_reg[106], loc_reg[107], loc_reg[108], loc_reg[109], loc_reg[110], loc_reg[111]} <= {loc_rdata[607:604], loc_rdata[603:600], loc_rdata[599:596], loc_rdata[595:592], loc_rdata[591:588], loc_rdata[587:584], loc_rdata[583:580], loc_rdata[579:576]};
        {loc_reg[112], loc_reg[113], loc_reg[114], loc_reg[115], loc_reg[116], loc_reg[117], loc_reg[118], loc_reg[119]} <= {loc_rdata[575:572], loc_rdata[571:568], loc_rdata[567:564], loc_rdata[563:560], loc_rdata[559:556], loc_rdata[555:552], loc_rdata[551:548], loc_rdata[547:544]};
        {loc_reg[120], loc_reg[121], loc_reg[122], loc_reg[123], loc_reg[124], loc_reg[125], loc_reg[126], loc_reg[127]} <= {loc_rdata[543:540], loc_rdata[539:536], loc_rdata[535:532], loc_rdata[531:528], loc_rdata[527:524], loc_rdata[523:520], loc_rdata[519:516], loc_rdata[515:512]};
        {loc_reg[128], loc_reg[129], loc_reg[130], loc_reg[131], loc_reg[132], loc_reg[133], loc_reg[134], loc_reg[135]} <= {loc_rdata[511:508], loc_rdata[507:504], loc_rdata[503:500], loc_rdata[499:496], loc_rdata[495:492], loc_rdata[491:488], loc_rdata[487:484], loc_rdata[483:480]};
        {loc_reg[136], loc_reg[137], loc_reg[138], loc_reg[139], loc_reg[140], loc_reg[141], loc_reg[142], loc_reg[143]} <= {loc_rdata[479:476], loc_rdata[475:472], loc_rdata[471:468], loc_rdata[467:464], loc_rdata[463:460], loc_rdata[459:456], loc_rdata[455:452], loc_rdata[451:448]};
        {loc_reg[144], loc_reg[145], loc_reg[146], loc_reg[147], loc_reg[148], loc_reg[149], loc_reg[150], loc_reg[151]} <= {loc_rdata[447:444], loc_rdata[443:440], loc_rdata[439:436], loc_rdata[435:432], loc_rdata[431:428], loc_rdata[427:424], loc_rdata[423:420], loc_rdata[419:416]};
        {loc_reg[152], loc_reg[153], loc_reg[154], loc_reg[155], loc_reg[156], loc_reg[157], loc_reg[158], loc_reg[159]} <= {loc_rdata[415:412], loc_rdata[411:408], loc_rdata[407:404], loc_rdata[403:400], loc_rdata[399:396], loc_rdata[395:392], loc_rdata[391:388], loc_rdata[387:384]};
        {loc_reg[160], loc_reg[161], loc_reg[162], loc_reg[163], loc_reg[164], loc_reg[165], loc_reg[166], loc_reg[167]} <= {loc_rdata[383:380], loc_rdata[379:376], loc_rdata[375:372], loc_rdata[371:368], loc_rdata[367:364], loc_rdata[363:360], loc_rdata[359:356], loc_rdata[355:352]};
        {loc_reg[168], loc_reg[169], loc_reg[170], loc_reg[171], loc_reg[172], loc_reg[173], loc_reg[174], loc_reg[175]} <= {loc_rdata[351:348], loc_rdata[347:344], loc_rdata[343:340], loc_rdata[339:336], loc_rdata[335:332], loc_rdata[331:328], loc_rdata[327:324], loc_rdata[323:320]};
        {loc_reg[176], loc_reg[177], loc_reg[178], loc_reg[179], loc_reg[180], loc_reg[181], loc_reg[182], loc_reg[183]} <= {loc_rdata[319:316], loc_rdata[315:312], loc_rdata[311:308], loc_rdata[307:304], loc_rdata[303:300], loc_rdata[299:296], loc_rdata[295:292], loc_rdata[291:288]};
        {loc_reg[184], loc_reg[185], loc_reg[186], loc_reg[187], loc_reg[188], loc_reg[189], loc_reg[190], loc_reg[191]} <= {loc_rdata[287:284], loc_rdata[283:280], loc_rdata[279:276], loc_rdata[275:272], loc_rdata[271:268], loc_rdata[267:264], loc_rdata[263:260], loc_rdata[259:256]};
        {loc_reg[192], loc_reg[193], loc_reg[194], loc_reg[195], loc_reg[196], loc_reg[197], loc_reg[198], loc_reg[199]} <= {loc_rdata[255:252], loc_rdata[251:248], loc_rdata[247:244], loc_rdata[243:240], loc_rdata[239:236], loc_rdata[235:232], loc_rdata[231:228], loc_rdata[227:224]};
        {loc_reg[200], loc_reg[201], loc_reg[202], loc_reg[203], loc_reg[204], loc_reg[205], loc_reg[206], loc_reg[207]} <= {loc_rdata[223:220], loc_rdata[219:216], loc_rdata[215:212], loc_rdata[211:208], loc_rdata[207:204], loc_rdata[203:200], loc_rdata[199:196], loc_rdata[195:192]};
        {loc_reg[208], loc_reg[209], loc_reg[210], loc_reg[211], loc_reg[212], loc_reg[213], loc_reg[214], loc_reg[215]} <= {loc_rdata[191:188], loc_rdata[187:184], loc_rdata[183:180], loc_rdata[179:176], loc_rdata[175:172], loc_rdata[171:168], loc_rdata[167:164], loc_rdata[163:160]};
        {loc_reg[216], loc_reg[217], loc_reg[218], loc_reg[219], loc_reg[220], loc_reg[221], loc_reg[222], loc_reg[223]} <= {loc_rdata[159:156], loc_rdata[155:152], loc_rdata[151:148], loc_rdata[147:144], loc_rdata[143:140], loc_rdata[139:136], loc_rdata[135:132], loc_rdata[131:128]};
        {loc_reg[224], loc_reg[225], loc_reg[226], loc_reg[227], loc_reg[228], loc_reg[229], loc_reg[230], loc_reg[231]} <= {loc_rdata[127:124], loc_rdata[123:120], loc_rdata[119:116], loc_rdata[115:112], loc_rdata[111:108], loc_rdata[107:104], loc_rdata[103:100], loc_rdata[99:96]};
        {loc_reg[232], loc_reg[233], loc_reg[234], loc_reg[235], loc_reg[236], loc_reg[237], loc_reg[238], loc_reg[239]} <= {loc_rdata[95:92], loc_rdata[91:88], loc_rdata[87:84], loc_rdata[83:80], loc_rdata[79:76], loc_rdata[75:72], loc_rdata[71:68], loc_rdata[67:64]};
        {loc_reg[240], loc_reg[241], loc_reg[242], loc_reg[243], loc_reg[244], loc_reg[245], loc_reg[246], loc_reg[247]} <= {loc_rdata[63:60], loc_rdata[59:56], loc_rdata[55:52], loc_rdata[51:48], loc_rdata[47:44], loc_rdata[43:40], loc_rdata[39:36], loc_rdata[35:32]};
        {loc_reg[248], loc_reg[249], loc_reg[250], loc_reg[251], loc_reg[252], loc_reg[253], loc_reg[254], loc_reg[255]} <= {loc_rdata[31:28], loc_rdata[27:24], loc_rdata[23:20], loc_rdata[19:16], loc_rdata[15:12], loc_rdata[11:8], loc_rdata[7:4], loc_rdata[3:0]};     
    end
end

// fsm
always@* begin
    case(state)
        IDLE: begin
            n_batch_finish = 0;
            n_ready = 0;
            if(en_in) begin
                n_state = DELAY1;
                n_sub_bat = 0;
            end else begin
                n_state = IDLE;
                n_sub_bat = 0;
            end
        end
		DELAY1: begin
			n_sub_bat = 0;
			n_batch_finish = 0;
			n_ready = 0;								
			n_state = SUB;
		end
        SUB: begin
            n_batch_finish = 0;
			n_ready = ((batch_num_reg > 0 && sub_bat == 1)) ? 1 : 0;
            n_state = (sub_bat == 15) ? DELAY2 : SUB;
			n_sub_bat = sub_bat + 1;
        end
		DELAY2: begin
			n_sub_bat = 0;
			n_batch_finish = 0;
			n_ready = 0;								
			n_state = CHECK;
		end
        CHECK: begin
          	n_sub_bat = 1;
			n_ready = 0;
            n_batch_finish = 0;
            n_state = (batch_num_reg == 8'd0) ? FIN : SUB;
        end
        FIN: begin
            n_sub_bat = sub_bat + 1;
            n_batch_finish = (sub_bat == 4'd4) ? 1 : 0;
            n_ready = (sub_bat == 4'd1) ? 1 : 0;
            n_state = (sub_bat == 4'd4) ? IDLE : FIN;
        end
        default: begin
            n_sub_bat = 0;
            n_batch_finish = 0;
            n_ready = 0;
            n_state = IDLE;
        end
    endcase
end

// COMB1: 256 X 16 to 1 mux so as to get n_loc_oh_reg
always@* begin
	case(loc_reg[0])
		4'd0: n_loc_oh_reg[0] = {15'd0, dist_reg[255]};
		4'd1: n_loc_oh_reg[0] = {14'd0, dist_reg[255], 1'd0};
		4'd2: n_loc_oh_reg[0] = {13'd0, dist_reg[255], 2'd0};
		4'd3: n_loc_oh_reg[0] = {12'd0, dist_reg[255], 3'd0};
		4'd4: n_loc_oh_reg[0] = {11'd0, dist_reg[255], 4'd0};
		4'd5: n_loc_oh_reg[0] = {10'd0, dist_reg[255], 5'd0};
		4'd6: n_loc_oh_reg[0] = {9'd0, dist_reg[255], 6'd0};
		4'd7: n_loc_oh_reg[0] = {8'd0, dist_reg[255], 7'd0};
		4'd8: n_loc_oh_reg[0] = {7'd0, dist_reg[255], 8'd0};
		4'd9: n_loc_oh_reg[0] = {6'd0, dist_reg[255], 9'd0};
		4'd10: n_loc_oh_reg[0] = {5'd0, dist_reg[255], 10'd0};
		4'd11: n_loc_oh_reg[0] = {4'd0, dist_reg[255], 11'd0};
		4'd12: n_loc_oh_reg[0] = {3'd0, dist_reg[255], 12'd0};
		4'd13: n_loc_oh_reg[0] = {2'd0, dist_reg[255], 13'd0};
		4'd14: n_loc_oh_reg[0] = {1'd0, dist_reg[255], 14'd0};
		4'd15: n_loc_oh_reg[0] = {dist_reg[255], 15'd0};
	endcase
	case(loc_reg[1])
		4'd0: n_loc_oh_reg[1] = {15'd0, dist_reg[254]};
		4'd1: n_loc_oh_reg[1] = {14'd0, dist_reg[254], 1'd0};
		4'd2: n_loc_oh_reg[1] = {13'd0, dist_reg[254], 2'd0};
		4'd3: n_loc_oh_reg[1] = {12'd0, dist_reg[254], 3'd0};
		4'd4: n_loc_oh_reg[1] = {11'd0, dist_reg[254], 4'd0};
		4'd5: n_loc_oh_reg[1] = {10'd0, dist_reg[254], 5'd0};
		4'd6: n_loc_oh_reg[1] = {9'd0, dist_reg[254], 6'd0};
		4'd7: n_loc_oh_reg[1] = {8'd0, dist_reg[254], 7'd0};
		4'd8: n_loc_oh_reg[1] = {7'd0, dist_reg[254], 8'd0};
		4'd9: n_loc_oh_reg[1] = {6'd0, dist_reg[254], 9'd0};
		4'd10: n_loc_oh_reg[1] = {5'd0, dist_reg[254], 10'd0};
		4'd11: n_loc_oh_reg[1] = {4'd0, dist_reg[254], 11'd0};
		4'd12: n_loc_oh_reg[1] = {3'd0, dist_reg[254], 12'd0};
		4'd13: n_loc_oh_reg[1] = {2'd0, dist_reg[254], 13'd0};
		4'd14: n_loc_oh_reg[1] = {1'd0, dist_reg[254], 14'd0};
		4'd15: n_loc_oh_reg[1] = {dist_reg[254], 15'd0};
	endcase
	case(loc_reg[2])
		4'd0: n_loc_oh_reg[2] = {15'd0, dist_reg[253]};
		4'd1: n_loc_oh_reg[2] = {14'd0, dist_reg[253], 1'd0};
		4'd2: n_loc_oh_reg[2] = {13'd0, dist_reg[253], 2'd0};
		4'd3: n_loc_oh_reg[2] = {12'd0, dist_reg[253], 3'd0};
		4'd4: n_loc_oh_reg[2] = {11'd0, dist_reg[253], 4'd0};
		4'd5: n_loc_oh_reg[2] = {10'd0, dist_reg[253], 5'd0};
		4'd6: n_loc_oh_reg[2] = {9'd0, dist_reg[253], 6'd0};
		4'd7: n_loc_oh_reg[2] = {8'd0, dist_reg[253], 7'd0};
		4'd8: n_loc_oh_reg[2] = {7'd0, dist_reg[253], 8'd0};
		4'd9: n_loc_oh_reg[2] = {6'd0, dist_reg[253], 9'd0};
		4'd10: n_loc_oh_reg[2] = {5'd0, dist_reg[253], 10'd0};
		4'd11: n_loc_oh_reg[2] = {4'd0, dist_reg[253], 11'd0};
		4'd12: n_loc_oh_reg[2] = {3'd0, dist_reg[253], 12'd0};
		4'd13: n_loc_oh_reg[2] = {2'd0, dist_reg[253], 13'd0};
		4'd14: n_loc_oh_reg[2] = {1'd0, dist_reg[253], 14'd0};
		4'd15: n_loc_oh_reg[2] = {dist_reg[253], 15'd0};
	endcase
	case(loc_reg[3])
		4'd0: n_loc_oh_reg[3] = {15'd0, dist_reg[252]};
		4'd1: n_loc_oh_reg[3] = {14'd0, dist_reg[252], 1'd0};
		4'd2: n_loc_oh_reg[3] = {13'd0, dist_reg[252], 2'd0};
		4'd3: n_loc_oh_reg[3] = {12'd0, dist_reg[252], 3'd0};
		4'd4: n_loc_oh_reg[3] = {11'd0, dist_reg[252], 4'd0};
		4'd5: n_loc_oh_reg[3] = {10'd0, dist_reg[252], 5'd0};
		4'd6: n_loc_oh_reg[3] = {9'd0, dist_reg[252], 6'd0};
		4'd7: n_loc_oh_reg[3] = {8'd0, dist_reg[252], 7'd0};
		4'd8: n_loc_oh_reg[3] = {7'd0, dist_reg[252], 8'd0};
		4'd9: n_loc_oh_reg[3] = {6'd0, dist_reg[252], 9'd0};
		4'd10: n_loc_oh_reg[3] = {5'd0, dist_reg[252], 10'd0};
		4'd11: n_loc_oh_reg[3] = {4'd0, dist_reg[252], 11'd0};
		4'd12: n_loc_oh_reg[3] = {3'd0, dist_reg[252], 12'd0};
		4'd13: n_loc_oh_reg[3] = {2'd0, dist_reg[252], 13'd0};
		4'd14: n_loc_oh_reg[3] = {1'd0, dist_reg[252], 14'd0};
		4'd15: n_loc_oh_reg[3] = {dist_reg[252], 15'd0};
	endcase
	case(loc_reg[4])
		4'd0: n_loc_oh_reg[4] = {15'd0, dist_reg[251]};
		4'd1: n_loc_oh_reg[4] = {14'd0, dist_reg[251], 1'd0};
		4'd2: n_loc_oh_reg[4] = {13'd0, dist_reg[251], 2'd0};
		4'd3: n_loc_oh_reg[4] = {12'd0, dist_reg[251], 3'd0};
		4'd4: n_loc_oh_reg[4] = {11'd0, dist_reg[251], 4'd0};
		4'd5: n_loc_oh_reg[4] = {10'd0, dist_reg[251], 5'd0};
		4'd6: n_loc_oh_reg[4] = {9'd0, dist_reg[251], 6'd0};
		4'd7: n_loc_oh_reg[4] = {8'd0, dist_reg[251], 7'd0};
		4'd8: n_loc_oh_reg[4] = {7'd0, dist_reg[251], 8'd0};
		4'd9: n_loc_oh_reg[4] = {6'd0, dist_reg[251], 9'd0};
		4'd10: n_loc_oh_reg[4] = {5'd0, dist_reg[251], 10'd0};
		4'd11: n_loc_oh_reg[4] = {4'd0, dist_reg[251], 11'd0};
		4'd12: n_loc_oh_reg[4] = {3'd0, dist_reg[251], 12'd0};
		4'd13: n_loc_oh_reg[4] = {2'd0, dist_reg[251], 13'd0};
		4'd14: n_loc_oh_reg[4] = {1'd0, dist_reg[251], 14'd0};
		4'd15: n_loc_oh_reg[4] = {dist_reg[251], 15'd0};
	endcase
	case(loc_reg[5])
		4'd0: n_loc_oh_reg[5] = {15'd0, dist_reg[250]};
		4'd1: n_loc_oh_reg[5] = {14'd0, dist_reg[250], 1'd0};
		4'd2: n_loc_oh_reg[5] = {13'd0, dist_reg[250], 2'd0};
		4'd3: n_loc_oh_reg[5] = {12'd0, dist_reg[250], 3'd0};
		4'd4: n_loc_oh_reg[5] = {11'd0, dist_reg[250], 4'd0};
		4'd5: n_loc_oh_reg[5] = {10'd0, dist_reg[250], 5'd0};
		4'd6: n_loc_oh_reg[5] = {9'd0, dist_reg[250], 6'd0};
		4'd7: n_loc_oh_reg[5] = {8'd0, dist_reg[250], 7'd0};
		4'd8: n_loc_oh_reg[5] = {7'd0, dist_reg[250], 8'd0};
		4'd9: n_loc_oh_reg[5] = {6'd0, dist_reg[250], 9'd0};
		4'd10: n_loc_oh_reg[5] = {5'd0, dist_reg[250], 10'd0};
		4'd11: n_loc_oh_reg[5] = {4'd0, dist_reg[250], 11'd0};
		4'd12: n_loc_oh_reg[5] = {3'd0, dist_reg[250], 12'd0};
		4'd13: n_loc_oh_reg[5] = {2'd0, dist_reg[250], 13'd0};
		4'd14: n_loc_oh_reg[5] = {1'd0, dist_reg[250], 14'd0};
		4'd15: n_loc_oh_reg[5] = {dist_reg[250], 15'd0};
	endcase
	case(loc_reg[6])
		4'd0: n_loc_oh_reg[6] = {15'd0, dist_reg[249]};
		4'd1: n_loc_oh_reg[6] = {14'd0, dist_reg[249], 1'd0};
		4'd2: n_loc_oh_reg[6] = {13'd0, dist_reg[249], 2'd0};
		4'd3: n_loc_oh_reg[6] = {12'd0, dist_reg[249], 3'd0};
		4'd4: n_loc_oh_reg[6] = {11'd0, dist_reg[249], 4'd0};
		4'd5: n_loc_oh_reg[6] = {10'd0, dist_reg[249], 5'd0};
		4'd6: n_loc_oh_reg[6] = {9'd0, dist_reg[249], 6'd0};
		4'd7: n_loc_oh_reg[6] = {8'd0, dist_reg[249], 7'd0};
		4'd8: n_loc_oh_reg[6] = {7'd0, dist_reg[249], 8'd0};
		4'd9: n_loc_oh_reg[6] = {6'd0, dist_reg[249], 9'd0};
		4'd10: n_loc_oh_reg[6] = {5'd0, dist_reg[249], 10'd0};
		4'd11: n_loc_oh_reg[6] = {4'd0, dist_reg[249], 11'd0};
		4'd12: n_loc_oh_reg[6] = {3'd0, dist_reg[249], 12'd0};
		4'd13: n_loc_oh_reg[6] = {2'd0, dist_reg[249], 13'd0};
		4'd14: n_loc_oh_reg[6] = {1'd0, dist_reg[249], 14'd0};
		4'd15: n_loc_oh_reg[6] = {dist_reg[249], 15'd0};
	endcase
	case(loc_reg[7])
		4'd0: n_loc_oh_reg[7] = {15'd0, dist_reg[248]};
		4'd1: n_loc_oh_reg[7] = {14'd0, dist_reg[248], 1'd0};
		4'd2: n_loc_oh_reg[7] = {13'd0, dist_reg[248], 2'd0};
		4'd3: n_loc_oh_reg[7] = {12'd0, dist_reg[248], 3'd0};
		4'd4: n_loc_oh_reg[7] = {11'd0, dist_reg[248], 4'd0};
		4'd5: n_loc_oh_reg[7] = {10'd0, dist_reg[248], 5'd0};
		4'd6: n_loc_oh_reg[7] = {9'd0, dist_reg[248], 6'd0};
		4'd7: n_loc_oh_reg[7] = {8'd0, dist_reg[248], 7'd0};
		4'd8: n_loc_oh_reg[7] = {7'd0, dist_reg[248], 8'd0};
		4'd9: n_loc_oh_reg[7] = {6'd0, dist_reg[248], 9'd0};
		4'd10: n_loc_oh_reg[7] = {5'd0, dist_reg[248], 10'd0};
		4'd11: n_loc_oh_reg[7] = {4'd0, dist_reg[248], 11'd0};
		4'd12: n_loc_oh_reg[7] = {3'd0, dist_reg[248], 12'd0};
		4'd13: n_loc_oh_reg[7] = {2'd0, dist_reg[248], 13'd0};
		4'd14: n_loc_oh_reg[7] = {1'd0, dist_reg[248], 14'd0};
		4'd15: n_loc_oh_reg[7] = {dist_reg[248], 15'd0};
	endcase
	case(loc_reg[8])
		4'd0: n_loc_oh_reg[8] = {15'd0, dist_reg[247]};
		4'd1: n_loc_oh_reg[8] = {14'd0, dist_reg[247], 1'd0};
		4'd2: n_loc_oh_reg[8] = {13'd0, dist_reg[247], 2'd0};
		4'd3: n_loc_oh_reg[8] = {12'd0, dist_reg[247], 3'd0};
		4'd4: n_loc_oh_reg[8] = {11'd0, dist_reg[247], 4'd0};
		4'd5: n_loc_oh_reg[8] = {10'd0, dist_reg[247], 5'd0};
		4'd6: n_loc_oh_reg[8] = {9'd0, dist_reg[247], 6'd0};
		4'd7: n_loc_oh_reg[8] = {8'd0, dist_reg[247], 7'd0};
		4'd8: n_loc_oh_reg[8] = {7'd0, dist_reg[247], 8'd0};
		4'd9: n_loc_oh_reg[8] = {6'd0, dist_reg[247], 9'd0};
		4'd10: n_loc_oh_reg[8] = {5'd0, dist_reg[247], 10'd0};
		4'd11: n_loc_oh_reg[8] = {4'd0, dist_reg[247], 11'd0};
		4'd12: n_loc_oh_reg[8] = {3'd0, dist_reg[247], 12'd0};
		4'd13: n_loc_oh_reg[8] = {2'd0, dist_reg[247], 13'd0};
		4'd14: n_loc_oh_reg[8] = {1'd0, dist_reg[247], 14'd0};
		4'd15: n_loc_oh_reg[8] = {dist_reg[247], 15'd0};
	endcase
	case(loc_reg[9])
		4'd0: n_loc_oh_reg[9] = {15'd0, dist_reg[246]};
		4'd1: n_loc_oh_reg[9] = {14'd0, dist_reg[246], 1'd0};
		4'd2: n_loc_oh_reg[9] = {13'd0, dist_reg[246], 2'd0};
		4'd3: n_loc_oh_reg[9] = {12'd0, dist_reg[246], 3'd0};
		4'd4: n_loc_oh_reg[9] = {11'd0, dist_reg[246], 4'd0};
		4'd5: n_loc_oh_reg[9] = {10'd0, dist_reg[246], 5'd0};
		4'd6: n_loc_oh_reg[9] = {9'd0, dist_reg[246], 6'd0};
		4'd7: n_loc_oh_reg[9] = {8'd0, dist_reg[246], 7'd0};
		4'd8: n_loc_oh_reg[9] = {7'd0, dist_reg[246], 8'd0};
		4'd9: n_loc_oh_reg[9] = {6'd0, dist_reg[246], 9'd0};
		4'd10: n_loc_oh_reg[9] = {5'd0, dist_reg[246], 10'd0};
		4'd11: n_loc_oh_reg[9] = {4'd0, dist_reg[246], 11'd0};
		4'd12: n_loc_oh_reg[9] = {3'd0, dist_reg[246], 12'd0};
		4'd13: n_loc_oh_reg[9] = {2'd0, dist_reg[246], 13'd0};
		4'd14: n_loc_oh_reg[9] = {1'd0, dist_reg[246], 14'd0};
		4'd15: n_loc_oh_reg[9] = {dist_reg[246], 15'd0};
	endcase
	case(loc_reg[10])
		4'd0: n_loc_oh_reg[10] = {15'd0, dist_reg[245]};
		4'd1: n_loc_oh_reg[10] = {14'd0, dist_reg[245], 1'd0};
		4'd2: n_loc_oh_reg[10] = {13'd0, dist_reg[245], 2'd0};
		4'd3: n_loc_oh_reg[10] = {12'd0, dist_reg[245], 3'd0};
		4'd4: n_loc_oh_reg[10] = {11'd0, dist_reg[245], 4'd0};
		4'd5: n_loc_oh_reg[10] = {10'd0, dist_reg[245], 5'd0};
		4'd6: n_loc_oh_reg[10] = {9'd0, dist_reg[245], 6'd0};
		4'd7: n_loc_oh_reg[10] = {8'd0, dist_reg[245], 7'd0};
		4'd8: n_loc_oh_reg[10] = {7'd0, dist_reg[245], 8'd0};
		4'd9: n_loc_oh_reg[10] = {6'd0, dist_reg[245], 9'd0};
		4'd10: n_loc_oh_reg[10] = {5'd0, dist_reg[245], 10'd0};
		4'd11: n_loc_oh_reg[10] = {4'd0, dist_reg[245], 11'd0};
		4'd12: n_loc_oh_reg[10] = {3'd0, dist_reg[245], 12'd0};
		4'd13: n_loc_oh_reg[10] = {2'd0, dist_reg[245], 13'd0};
		4'd14: n_loc_oh_reg[10] = {1'd0, dist_reg[245], 14'd0};
		4'd15: n_loc_oh_reg[10] = {dist_reg[245], 15'd0};
	endcase
	case(loc_reg[11])
		4'd0: n_loc_oh_reg[11] = {15'd0, dist_reg[244]};
		4'd1: n_loc_oh_reg[11] = {14'd0, dist_reg[244], 1'd0};
		4'd2: n_loc_oh_reg[11] = {13'd0, dist_reg[244], 2'd0};
		4'd3: n_loc_oh_reg[11] = {12'd0, dist_reg[244], 3'd0};
		4'd4: n_loc_oh_reg[11] = {11'd0, dist_reg[244], 4'd0};
		4'd5: n_loc_oh_reg[11] = {10'd0, dist_reg[244], 5'd0};
		4'd6: n_loc_oh_reg[11] = {9'd0, dist_reg[244], 6'd0};
		4'd7: n_loc_oh_reg[11] = {8'd0, dist_reg[244], 7'd0};
		4'd8: n_loc_oh_reg[11] = {7'd0, dist_reg[244], 8'd0};
		4'd9: n_loc_oh_reg[11] = {6'd0, dist_reg[244], 9'd0};
		4'd10: n_loc_oh_reg[11] = {5'd0, dist_reg[244], 10'd0};
		4'd11: n_loc_oh_reg[11] = {4'd0, dist_reg[244], 11'd0};
		4'd12: n_loc_oh_reg[11] = {3'd0, dist_reg[244], 12'd0};
		4'd13: n_loc_oh_reg[11] = {2'd0, dist_reg[244], 13'd0};
		4'd14: n_loc_oh_reg[11] = {1'd0, dist_reg[244], 14'd0};
		4'd15: n_loc_oh_reg[11] = {dist_reg[244], 15'd0};
	endcase
	case(loc_reg[12])
		4'd0: n_loc_oh_reg[12] = {15'd0, dist_reg[243]};
		4'd1: n_loc_oh_reg[12] = {14'd0, dist_reg[243], 1'd0};
		4'd2: n_loc_oh_reg[12] = {13'd0, dist_reg[243], 2'd0};
		4'd3: n_loc_oh_reg[12] = {12'd0, dist_reg[243], 3'd0};
		4'd4: n_loc_oh_reg[12] = {11'd0, dist_reg[243], 4'd0};
		4'd5: n_loc_oh_reg[12] = {10'd0, dist_reg[243], 5'd0};
		4'd6: n_loc_oh_reg[12] = {9'd0, dist_reg[243], 6'd0};
		4'd7: n_loc_oh_reg[12] = {8'd0, dist_reg[243], 7'd0};
		4'd8: n_loc_oh_reg[12] = {7'd0, dist_reg[243], 8'd0};
		4'd9: n_loc_oh_reg[12] = {6'd0, dist_reg[243], 9'd0};
		4'd10: n_loc_oh_reg[12] = {5'd0, dist_reg[243], 10'd0};
		4'd11: n_loc_oh_reg[12] = {4'd0, dist_reg[243], 11'd0};
		4'd12: n_loc_oh_reg[12] = {3'd0, dist_reg[243], 12'd0};
		4'd13: n_loc_oh_reg[12] = {2'd0, dist_reg[243], 13'd0};
		4'd14: n_loc_oh_reg[12] = {1'd0, dist_reg[243], 14'd0};
		4'd15: n_loc_oh_reg[12] = {dist_reg[243], 15'd0};
	endcase
	case(loc_reg[13])
		4'd0: n_loc_oh_reg[13] = {15'd0, dist_reg[242]};
		4'd1: n_loc_oh_reg[13] = {14'd0, dist_reg[242], 1'd0};
		4'd2: n_loc_oh_reg[13] = {13'd0, dist_reg[242], 2'd0};
		4'd3: n_loc_oh_reg[13] = {12'd0, dist_reg[242], 3'd0};
		4'd4: n_loc_oh_reg[13] = {11'd0, dist_reg[242], 4'd0};
		4'd5: n_loc_oh_reg[13] = {10'd0, dist_reg[242], 5'd0};
		4'd6: n_loc_oh_reg[13] = {9'd0, dist_reg[242], 6'd0};
		4'd7: n_loc_oh_reg[13] = {8'd0, dist_reg[242], 7'd0};
		4'd8: n_loc_oh_reg[13] = {7'd0, dist_reg[242], 8'd0};
		4'd9: n_loc_oh_reg[13] = {6'd0, dist_reg[242], 9'd0};
		4'd10: n_loc_oh_reg[13] = {5'd0, dist_reg[242], 10'd0};
		4'd11: n_loc_oh_reg[13] = {4'd0, dist_reg[242], 11'd0};
		4'd12: n_loc_oh_reg[13] = {3'd0, dist_reg[242], 12'd0};
		4'd13: n_loc_oh_reg[13] = {2'd0, dist_reg[242], 13'd0};
		4'd14: n_loc_oh_reg[13] = {1'd0, dist_reg[242], 14'd0};
		4'd15: n_loc_oh_reg[13] = {dist_reg[242], 15'd0};
	endcase
	case(loc_reg[14])
		4'd0: n_loc_oh_reg[14] = {15'd0, dist_reg[241]};
		4'd1: n_loc_oh_reg[14] = {14'd0, dist_reg[241], 1'd0};
		4'd2: n_loc_oh_reg[14] = {13'd0, dist_reg[241], 2'd0};
		4'd3: n_loc_oh_reg[14] = {12'd0, dist_reg[241], 3'd0};
		4'd4: n_loc_oh_reg[14] = {11'd0, dist_reg[241], 4'd0};
		4'd5: n_loc_oh_reg[14] = {10'd0, dist_reg[241], 5'd0};
		4'd6: n_loc_oh_reg[14] = {9'd0, dist_reg[241], 6'd0};
		4'd7: n_loc_oh_reg[14] = {8'd0, dist_reg[241], 7'd0};
		4'd8: n_loc_oh_reg[14] = {7'd0, dist_reg[241], 8'd0};
		4'd9: n_loc_oh_reg[14] = {6'd0, dist_reg[241], 9'd0};
		4'd10: n_loc_oh_reg[14] = {5'd0, dist_reg[241], 10'd0};
		4'd11: n_loc_oh_reg[14] = {4'd0, dist_reg[241], 11'd0};
		4'd12: n_loc_oh_reg[14] = {3'd0, dist_reg[241], 12'd0};
		4'd13: n_loc_oh_reg[14] = {2'd0, dist_reg[241], 13'd0};
		4'd14: n_loc_oh_reg[14] = {1'd0, dist_reg[241], 14'd0};
		4'd15: n_loc_oh_reg[14] = {dist_reg[241], 15'd0};
	endcase
	case(loc_reg[15])
		4'd0: n_loc_oh_reg[15] = {15'd0, dist_reg[240]};
		4'd1: n_loc_oh_reg[15] = {14'd0, dist_reg[240], 1'd0};
		4'd2: n_loc_oh_reg[15] = {13'd0, dist_reg[240], 2'd0};
		4'd3: n_loc_oh_reg[15] = {12'd0, dist_reg[240], 3'd0};
		4'd4: n_loc_oh_reg[15] = {11'd0, dist_reg[240], 4'd0};
		4'd5: n_loc_oh_reg[15] = {10'd0, dist_reg[240], 5'd0};
		4'd6: n_loc_oh_reg[15] = {9'd0, dist_reg[240], 6'd0};
		4'd7: n_loc_oh_reg[15] = {8'd0, dist_reg[240], 7'd0};
		4'd8: n_loc_oh_reg[15] = {7'd0, dist_reg[240], 8'd0};
		4'd9: n_loc_oh_reg[15] = {6'd0, dist_reg[240], 9'd0};
		4'd10: n_loc_oh_reg[15] = {5'd0, dist_reg[240], 10'd0};
		4'd11: n_loc_oh_reg[15] = {4'd0, dist_reg[240], 11'd0};
		4'd12: n_loc_oh_reg[15] = {3'd0, dist_reg[240], 12'd0};
		4'd13: n_loc_oh_reg[15] = {2'd0, dist_reg[240], 13'd0};
		4'd14: n_loc_oh_reg[15] = {1'd0, dist_reg[240], 14'd0};
		4'd15: n_loc_oh_reg[15] = {dist_reg[240], 15'd0};
	endcase
	case(loc_reg[16])
		4'd0: n_loc_oh_reg[16] = {15'd0, dist_reg[239]};
		4'd1: n_loc_oh_reg[16] = {14'd0, dist_reg[239], 1'd0};
		4'd2: n_loc_oh_reg[16] = {13'd0, dist_reg[239], 2'd0};
		4'd3: n_loc_oh_reg[16] = {12'd0, dist_reg[239], 3'd0};
		4'd4: n_loc_oh_reg[16] = {11'd0, dist_reg[239], 4'd0};
		4'd5: n_loc_oh_reg[16] = {10'd0, dist_reg[239], 5'd0};
		4'd6: n_loc_oh_reg[16] = {9'd0, dist_reg[239], 6'd0};
		4'd7: n_loc_oh_reg[16] = {8'd0, dist_reg[239], 7'd0};
		4'd8: n_loc_oh_reg[16] = {7'd0, dist_reg[239], 8'd0};
		4'd9: n_loc_oh_reg[16] = {6'd0, dist_reg[239], 9'd0};
		4'd10: n_loc_oh_reg[16] = {5'd0, dist_reg[239], 10'd0};
		4'd11: n_loc_oh_reg[16] = {4'd0, dist_reg[239], 11'd0};
		4'd12: n_loc_oh_reg[16] = {3'd0, dist_reg[239], 12'd0};
		4'd13: n_loc_oh_reg[16] = {2'd0, dist_reg[239], 13'd0};
		4'd14: n_loc_oh_reg[16] = {1'd0, dist_reg[239], 14'd0};
		4'd15: n_loc_oh_reg[16] = {dist_reg[239], 15'd0};
	endcase
	case(loc_reg[17])
		4'd0: n_loc_oh_reg[17] = {15'd0, dist_reg[238]};
		4'd1: n_loc_oh_reg[17] = {14'd0, dist_reg[238], 1'd0};
		4'd2: n_loc_oh_reg[17] = {13'd0, dist_reg[238], 2'd0};
		4'd3: n_loc_oh_reg[17] = {12'd0, dist_reg[238], 3'd0};
		4'd4: n_loc_oh_reg[17] = {11'd0, dist_reg[238], 4'd0};
		4'd5: n_loc_oh_reg[17] = {10'd0, dist_reg[238], 5'd0};
		4'd6: n_loc_oh_reg[17] = {9'd0, dist_reg[238], 6'd0};
		4'd7: n_loc_oh_reg[17] = {8'd0, dist_reg[238], 7'd0};
		4'd8: n_loc_oh_reg[17] = {7'd0, dist_reg[238], 8'd0};
		4'd9: n_loc_oh_reg[17] = {6'd0, dist_reg[238], 9'd0};
		4'd10: n_loc_oh_reg[17] = {5'd0, dist_reg[238], 10'd0};
		4'd11: n_loc_oh_reg[17] = {4'd0, dist_reg[238], 11'd0};
		4'd12: n_loc_oh_reg[17] = {3'd0, dist_reg[238], 12'd0};
		4'd13: n_loc_oh_reg[17] = {2'd0, dist_reg[238], 13'd0};
		4'd14: n_loc_oh_reg[17] = {1'd0, dist_reg[238], 14'd0};
		4'd15: n_loc_oh_reg[17] = {dist_reg[238], 15'd0};
	endcase
	case(loc_reg[18])
		4'd0: n_loc_oh_reg[18] = {15'd0, dist_reg[237]};
		4'd1: n_loc_oh_reg[18] = {14'd0, dist_reg[237], 1'd0};
		4'd2: n_loc_oh_reg[18] = {13'd0, dist_reg[237], 2'd0};
		4'd3: n_loc_oh_reg[18] = {12'd0, dist_reg[237], 3'd0};
		4'd4: n_loc_oh_reg[18] = {11'd0, dist_reg[237], 4'd0};
		4'd5: n_loc_oh_reg[18] = {10'd0, dist_reg[237], 5'd0};
		4'd6: n_loc_oh_reg[18] = {9'd0, dist_reg[237], 6'd0};
		4'd7: n_loc_oh_reg[18] = {8'd0, dist_reg[237], 7'd0};
		4'd8: n_loc_oh_reg[18] = {7'd0, dist_reg[237], 8'd0};
		4'd9: n_loc_oh_reg[18] = {6'd0, dist_reg[237], 9'd0};
		4'd10: n_loc_oh_reg[18] = {5'd0, dist_reg[237], 10'd0};
		4'd11: n_loc_oh_reg[18] = {4'd0, dist_reg[237], 11'd0};
		4'd12: n_loc_oh_reg[18] = {3'd0, dist_reg[237], 12'd0};
		4'd13: n_loc_oh_reg[18] = {2'd0, dist_reg[237], 13'd0};
		4'd14: n_loc_oh_reg[18] = {1'd0, dist_reg[237], 14'd0};
		4'd15: n_loc_oh_reg[18] = {dist_reg[237], 15'd0};
	endcase
	case(loc_reg[19])
		4'd0: n_loc_oh_reg[19] = {15'd0, dist_reg[236]};
		4'd1: n_loc_oh_reg[19] = {14'd0, dist_reg[236], 1'd0};
		4'd2: n_loc_oh_reg[19] = {13'd0, dist_reg[236], 2'd0};
		4'd3: n_loc_oh_reg[19] = {12'd0, dist_reg[236], 3'd0};
		4'd4: n_loc_oh_reg[19] = {11'd0, dist_reg[236], 4'd0};
		4'd5: n_loc_oh_reg[19] = {10'd0, dist_reg[236], 5'd0};
		4'd6: n_loc_oh_reg[19] = {9'd0, dist_reg[236], 6'd0};
		4'd7: n_loc_oh_reg[19] = {8'd0, dist_reg[236], 7'd0};
		4'd8: n_loc_oh_reg[19] = {7'd0, dist_reg[236], 8'd0};
		4'd9: n_loc_oh_reg[19] = {6'd0, dist_reg[236], 9'd0};
		4'd10: n_loc_oh_reg[19] = {5'd0, dist_reg[236], 10'd0};
		4'd11: n_loc_oh_reg[19] = {4'd0, dist_reg[236], 11'd0};
		4'd12: n_loc_oh_reg[19] = {3'd0, dist_reg[236], 12'd0};
		4'd13: n_loc_oh_reg[19] = {2'd0, dist_reg[236], 13'd0};
		4'd14: n_loc_oh_reg[19] = {1'd0, dist_reg[236], 14'd0};
		4'd15: n_loc_oh_reg[19] = {dist_reg[236], 15'd0};
	endcase
	case(loc_reg[20])
		4'd0: n_loc_oh_reg[20] = {15'd0, dist_reg[235]};
		4'd1: n_loc_oh_reg[20] = {14'd0, dist_reg[235], 1'd0};
		4'd2: n_loc_oh_reg[20] = {13'd0, dist_reg[235], 2'd0};
		4'd3: n_loc_oh_reg[20] = {12'd0, dist_reg[235], 3'd0};
		4'd4: n_loc_oh_reg[20] = {11'd0, dist_reg[235], 4'd0};
		4'd5: n_loc_oh_reg[20] = {10'd0, dist_reg[235], 5'd0};
		4'd6: n_loc_oh_reg[20] = {9'd0, dist_reg[235], 6'd0};
		4'd7: n_loc_oh_reg[20] = {8'd0, dist_reg[235], 7'd0};
		4'd8: n_loc_oh_reg[20] = {7'd0, dist_reg[235], 8'd0};
		4'd9: n_loc_oh_reg[20] = {6'd0, dist_reg[235], 9'd0};
		4'd10: n_loc_oh_reg[20] = {5'd0, dist_reg[235], 10'd0};
		4'd11: n_loc_oh_reg[20] = {4'd0, dist_reg[235], 11'd0};
		4'd12: n_loc_oh_reg[20] = {3'd0, dist_reg[235], 12'd0};
		4'd13: n_loc_oh_reg[20] = {2'd0, dist_reg[235], 13'd0};
		4'd14: n_loc_oh_reg[20] = {1'd0, dist_reg[235], 14'd0};
		4'd15: n_loc_oh_reg[20] = {dist_reg[235], 15'd0};
	endcase
	case(loc_reg[21])
		4'd0: n_loc_oh_reg[21] = {15'd0, dist_reg[234]};
		4'd1: n_loc_oh_reg[21] = {14'd0, dist_reg[234], 1'd0};
		4'd2: n_loc_oh_reg[21] = {13'd0, dist_reg[234], 2'd0};
		4'd3: n_loc_oh_reg[21] = {12'd0, dist_reg[234], 3'd0};
		4'd4: n_loc_oh_reg[21] = {11'd0, dist_reg[234], 4'd0};
		4'd5: n_loc_oh_reg[21] = {10'd0, dist_reg[234], 5'd0};
		4'd6: n_loc_oh_reg[21] = {9'd0, dist_reg[234], 6'd0};
		4'd7: n_loc_oh_reg[21] = {8'd0, dist_reg[234], 7'd0};
		4'd8: n_loc_oh_reg[21] = {7'd0, dist_reg[234], 8'd0};
		4'd9: n_loc_oh_reg[21] = {6'd0, dist_reg[234], 9'd0};
		4'd10: n_loc_oh_reg[21] = {5'd0, dist_reg[234], 10'd0};
		4'd11: n_loc_oh_reg[21] = {4'd0, dist_reg[234], 11'd0};
		4'd12: n_loc_oh_reg[21] = {3'd0, dist_reg[234], 12'd0};
		4'd13: n_loc_oh_reg[21] = {2'd0, dist_reg[234], 13'd0};
		4'd14: n_loc_oh_reg[21] = {1'd0, dist_reg[234], 14'd0};
		4'd15: n_loc_oh_reg[21] = {dist_reg[234], 15'd0};
	endcase
	case(loc_reg[22])
		4'd0: n_loc_oh_reg[22] = {15'd0, dist_reg[233]};
		4'd1: n_loc_oh_reg[22] = {14'd0, dist_reg[233], 1'd0};
		4'd2: n_loc_oh_reg[22] = {13'd0, dist_reg[233], 2'd0};
		4'd3: n_loc_oh_reg[22] = {12'd0, dist_reg[233], 3'd0};
		4'd4: n_loc_oh_reg[22] = {11'd0, dist_reg[233], 4'd0};
		4'd5: n_loc_oh_reg[22] = {10'd0, dist_reg[233], 5'd0};
		4'd6: n_loc_oh_reg[22] = {9'd0, dist_reg[233], 6'd0};
		4'd7: n_loc_oh_reg[22] = {8'd0, dist_reg[233], 7'd0};
		4'd8: n_loc_oh_reg[22] = {7'd0, dist_reg[233], 8'd0};
		4'd9: n_loc_oh_reg[22] = {6'd0, dist_reg[233], 9'd0};
		4'd10: n_loc_oh_reg[22] = {5'd0, dist_reg[233], 10'd0};
		4'd11: n_loc_oh_reg[22] = {4'd0, dist_reg[233], 11'd0};
		4'd12: n_loc_oh_reg[22] = {3'd0, dist_reg[233], 12'd0};
		4'd13: n_loc_oh_reg[22] = {2'd0, dist_reg[233], 13'd0};
		4'd14: n_loc_oh_reg[22] = {1'd0, dist_reg[233], 14'd0};
		4'd15: n_loc_oh_reg[22] = {dist_reg[233], 15'd0};
	endcase
	case(loc_reg[23])
		4'd0: n_loc_oh_reg[23] = {15'd0, dist_reg[232]};
		4'd1: n_loc_oh_reg[23] = {14'd0, dist_reg[232], 1'd0};
		4'd2: n_loc_oh_reg[23] = {13'd0, dist_reg[232], 2'd0};
		4'd3: n_loc_oh_reg[23] = {12'd0, dist_reg[232], 3'd0};
		4'd4: n_loc_oh_reg[23] = {11'd0, dist_reg[232], 4'd0};
		4'd5: n_loc_oh_reg[23] = {10'd0, dist_reg[232], 5'd0};
		4'd6: n_loc_oh_reg[23] = {9'd0, dist_reg[232], 6'd0};
		4'd7: n_loc_oh_reg[23] = {8'd0, dist_reg[232], 7'd0};
		4'd8: n_loc_oh_reg[23] = {7'd0, dist_reg[232], 8'd0};
		4'd9: n_loc_oh_reg[23] = {6'd0, dist_reg[232], 9'd0};
		4'd10: n_loc_oh_reg[23] = {5'd0, dist_reg[232], 10'd0};
		4'd11: n_loc_oh_reg[23] = {4'd0, dist_reg[232], 11'd0};
		4'd12: n_loc_oh_reg[23] = {3'd0, dist_reg[232], 12'd0};
		4'd13: n_loc_oh_reg[23] = {2'd0, dist_reg[232], 13'd0};
		4'd14: n_loc_oh_reg[23] = {1'd0, dist_reg[232], 14'd0};
		4'd15: n_loc_oh_reg[23] = {dist_reg[232], 15'd0};
	endcase
	case(loc_reg[24])
		4'd0: n_loc_oh_reg[24] = {15'd0, dist_reg[231]};
		4'd1: n_loc_oh_reg[24] = {14'd0, dist_reg[231], 1'd0};
		4'd2: n_loc_oh_reg[24] = {13'd0, dist_reg[231], 2'd0};
		4'd3: n_loc_oh_reg[24] = {12'd0, dist_reg[231], 3'd0};
		4'd4: n_loc_oh_reg[24] = {11'd0, dist_reg[231], 4'd0};
		4'd5: n_loc_oh_reg[24] = {10'd0, dist_reg[231], 5'd0};
		4'd6: n_loc_oh_reg[24] = {9'd0, dist_reg[231], 6'd0};
		4'd7: n_loc_oh_reg[24] = {8'd0, dist_reg[231], 7'd0};
		4'd8: n_loc_oh_reg[24] = {7'd0, dist_reg[231], 8'd0};
		4'd9: n_loc_oh_reg[24] = {6'd0, dist_reg[231], 9'd0};
		4'd10: n_loc_oh_reg[24] = {5'd0, dist_reg[231], 10'd0};
		4'd11: n_loc_oh_reg[24] = {4'd0, dist_reg[231], 11'd0};
		4'd12: n_loc_oh_reg[24] = {3'd0, dist_reg[231], 12'd0};
		4'd13: n_loc_oh_reg[24] = {2'd0, dist_reg[231], 13'd0};
		4'd14: n_loc_oh_reg[24] = {1'd0, dist_reg[231], 14'd0};
		4'd15: n_loc_oh_reg[24] = {dist_reg[231], 15'd0};
	endcase
	case(loc_reg[25])
		4'd0: n_loc_oh_reg[25] = {15'd0, dist_reg[230]};
		4'd1: n_loc_oh_reg[25] = {14'd0, dist_reg[230], 1'd0};
		4'd2: n_loc_oh_reg[25] = {13'd0, dist_reg[230], 2'd0};
		4'd3: n_loc_oh_reg[25] = {12'd0, dist_reg[230], 3'd0};
		4'd4: n_loc_oh_reg[25] = {11'd0, dist_reg[230], 4'd0};
		4'd5: n_loc_oh_reg[25] = {10'd0, dist_reg[230], 5'd0};
		4'd6: n_loc_oh_reg[25] = {9'd0, dist_reg[230], 6'd0};
		4'd7: n_loc_oh_reg[25] = {8'd0, dist_reg[230], 7'd0};
		4'd8: n_loc_oh_reg[25] = {7'd0, dist_reg[230], 8'd0};
		4'd9: n_loc_oh_reg[25] = {6'd0, dist_reg[230], 9'd0};
		4'd10: n_loc_oh_reg[25] = {5'd0, dist_reg[230], 10'd0};
		4'd11: n_loc_oh_reg[25] = {4'd0, dist_reg[230], 11'd0};
		4'd12: n_loc_oh_reg[25] = {3'd0, dist_reg[230], 12'd0};
		4'd13: n_loc_oh_reg[25] = {2'd0, dist_reg[230], 13'd0};
		4'd14: n_loc_oh_reg[25] = {1'd0, dist_reg[230], 14'd0};
		4'd15: n_loc_oh_reg[25] = {dist_reg[230], 15'd0};
	endcase
	case(loc_reg[26])
		4'd0: n_loc_oh_reg[26] = {15'd0, dist_reg[229]};
		4'd1: n_loc_oh_reg[26] = {14'd0, dist_reg[229], 1'd0};
		4'd2: n_loc_oh_reg[26] = {13'd0, dist_reg[229], 2'd0};
		4'd3: n_loc_oh_reg[26] = {12'd0, dist_reg[229], 3'd0};
		4'd4: n_loc_oh_reg[26] = {11'd0, dist_reg[229], 4'd0};
		4'd5: n_loc_oh_reg[26] = {10'd0, dist_reg[229], 5'd0};
		4'd6: n_loc_oh_reg[26] = {9'd0, dist_reg[229], 6'd0};
		4'd7: n_loc_oh_reg[26] = {8'd0, dist_reg[229], 7'd0};
		4'd8: n_loc_oh_reg[26] = {7'd0, dist_reg[229], 8'd0};
		4'd9: n_loc_oh_reg[26] = {6'd0, dist_reg[229], 9'd0};
		4'd10: n_loc_oh_reg[26] = {5'd0, dist_reg[229], 10'd0};
		4'd11: n_loc_oh_reg[26] = {4'd0, dist_reg[229], 11'd0};
		4'd12: n_loc_oh_reg[26] = {3'd0, dist_reg[229], 12'd0};
		4'd13: n_loc_oh_reg[26] = {2'd0, dist_reg[229], 13'd0};
		4'd14: n_loc_oh_reg[26] = {1'd0, dist_reg[229], 14'd0};
		4'd15: n_loc_oh_reg[26] = {dist_reg[229], 15'd0};
	endcase
	case(loc_reg[27])
		4'd0: n_loc_oh_reg[27] = {15'd0, dist_reg[228]};
		4'd1: n_loc_oh_reg[27] = {14'd0, dist_reg[228], 1'd0};
		4'd2: n_loc_oh_reg[27] = {13'd0, dist_reg[228], 2'd0};
		4'd3: n_loc_oh_reg[27] = {12'd0, dist_reg[228], 3'd0};
		4'd4: n_loc_oh_reg[27] = {11'd0, dist_reg[228], 4'd0};
		4'd5: n_loc_oh_reg[27] = {10'd0, dist_reg[228], 5'd0};
		4'd6: n_loc_oh_reg[27] = {9'd0, dist_reg[228], 6'd0};
		4'd7: n_loc_oh_reg[27] = {8'd0, dist_reg[228], 7'd0};
		4'd8: n_loc_oh_reg[27] = {7'd0, dist_reg[228], 8'd0};
		4'd9: n_loc_oh_reg[27] = {6'd0, dist_reg[228], 9'd0};
		4'd10: n_loc_oh_reg[27] = {5'd0, dist_reg[228], 10'd0};
		4'd11: n_loc_oh_reg[27] = {4'd0, dist_reg[228], 11'd0};
		4'd12: n_loc_oh_reg[27] = {3'd0, dist_reg[228], 12'd0};
		4'd13: n_loc_oh_reg[27] = {2'd0, dist_reg[228], 13'd0};
		4'd14: n_loc_oh_reg[27] = {1'd0, dist_reg[228], 14'd0};
		4'd15: n_loc_oh_reg[27] = {dist_reg[228], 15'd0};
	endcase
	case(loc_reg[28])
		4'd0: n_loc_oh_reg[28] = {15'd0, dist_reg[227]};
		4'd1: n_loc_oh_reg[28] = {14'd0, dist_reg[227], 1'd0};
		4'd2: n_loc_oh_reg[28] = {13'd0, dist_reg[227], 2'd0};
		4'd3: n_loc_oh_reg[28] = {12'd0, dist_reg[227], 3'd0};
		4'd4: n_loc_oh_reg[28] = {11'd0, dist_reg[227], 4'd0};
		4'd5: n_loc_oh_reg[28] = {10'd0, dist_reg[227], 5'd0};
		4'd6: n_loc_oh_reg[28] = {9'd0, dist_reg[227], 6'd0};
		4'd7: n_loc_oh_reg[28] = {8'd0, dist_reg[227], 7'd0};
		4'd8: n_loc_oh_reg[28] = {7'd0, dist_reg[227], 8'd0};
		4'd9: n_loc_oh_reg[28] = {6'd0, dist_reg[227], 9'd0};
		4'd10: n_loc_oh_reg[28] = {5'd0, dist_reg[227], 10'd0};
		4'd11: n_loc_oh_reg[28] = {4'd0, dist_reg[227], 11'd0};
		4'd12: n_loc_oh_reg[28] = {3'd0, dist_reg[227], 12'd0};
		4'd13: n_loc_oh_reg[28] = {2'd0, dist_reg[227], 13'd0};
		4'd14: n_loc_oh_reg[28] = {1'd0, dist_reg[227], 14'd0};
		4'd15: n_loc_oh_reg[28] = {dist_reg[227], 15'd0};
	endcase
	case(loc_reg[29])
		4'd0: n_loc_oh_reg[29] = {15'd0, dist_reg[226]};
		4'd1: n_loc_oh_reg[29] = {14'd0, dist_reg[226], 1'd0};
		4'd2: n_loc_oh_reg[29] = {13'd0, dist_reg[226], 2'd0};
		4'd3: n_loc_oh_reg[29] = {12'd0, dist_reg[226], 3'd0};
		4'd4: n_loc_oh_reg[29] = {11'd0, dist_reg[226], 4'd0};
		4'd5: n_loc_oh_reg[29] = {10'd0, dist_reg[226], 5'd0};
		4'd6: n_loc_oh_reg[29] = {9'd0, dist_reg[226], 6'd0};
		4'd7: n_loc_oh_reg[29] = {8'd0, dist_reg[226], 7'd0};
		4'd8: n_loc_oh_reg[29] = {7'd0, dist_reg[226], 8'd0};
		4'd9: n_loc_oh_reg[29] = {6'd0, dist_reg[226], 9'd0};
		4'd10: n_loc_oh_reg[29] = {5'd0, dist_reg[226], 10'd0};
		4'd11: n_loc_oh_reg[29] = {4'd0, dist_reg[226], 11'd0};
		4'd12: n_loc_oh_reg[29] = {3'd0, dist_reg[226], 12'd0};
		4'd13: n_loc_oh_reg[29] = {2'd0, dist_reg[226], 13'd0};
		4'd14: n_loc_oh_reg[29] = {1'd0, dist_reg[226], 14'd0};
		4'd15: n_loc_oh_reg[29] = {dist_reg[226], 15'd0};
	endcase
	case(loc_reg[30])
		4'd0: n_loc_oh_reg[30] = {15'd0, dist_reg[225]};
		4'd1: n_loc_oh_reg[30] = {14'd0, dist_reg[225], 1'd0};
		4'd2: n_loc_oh_reg[30] = {13'd0, dist_reg[225], 2'd0};
		4'd3: n_loc_oh_reg[30] = {12'd0, dist_reg[225], 3'd0};
		4'd4: n_loc_oh_reg[30] = {11'd0, dist_reg[225], 4'd0};
		4'd5: n_loc_oh_reg[30] = {10'd0, dist_reg[225], 5'd0};
		4'd6: n_loc_oh_reg[30] = {9'd0, dist_reg[225], 6'd0};
		4'd7: n_loc_oh_reg[30] = {8'd0, dist_reg[225], 7'd0};
		4'd8: n_loc_oh_reg[30] = {7'd0, dist_reg[225], 8'd0};
		4'd9: n_loc_oh_reg[30] = {6'd0, dist_reg[225], 9'd0};
		4'd10: n_loc_oh_reg[30] = {5'd0, dist_reg[225], 10'd0};
		4'd11: n_loc_oh_reg[30] = {4'd0, dist_reg[225], 11'd0};
		4'd12: n_loc_oh_reg[30] = {3'd0, dist_reg[225], 12'd0};
		4'd13: n_loc_oh_reg[30] = {2'd0, dist_reg[225], 13'd0};
		4'd14: n_loc_oh_reg[30] = {1'd0, dist_reg[225], 14'd0};
		4'd15: n_loc_oh_reg[30] = {dist_reg[225], 15'd0};
	endcase
	case(loc_reg[31])
		4'd0: n_loc_oh_reg[31] = {15'd0, dist_reg[224]};
		4'd1: n_loc_oh_reg[31] = {14'd0, dist_reg[224], 1'd0};
		4'd2: n_loc_oh_reg[31] = {13'd0, dist_reg[224], 2'd0};
		4'd3: n_loc_oh_reg[31] = {12'd0, dist_reg[224], 3'd0};
		4'd4: n_loc_oh_reg[31] = {11'd0, dist_reg[224], 4'd0};
		4'd5: n_loc_oh_reg[31] = {10'd0, dist_reg[224], 5'd0};
		4'd6: n_loc_oh_reg[31] = {9'd0, dist_reg[224], 6'd0};
		4'd7: n_loc_oh_reg[31] = {8'd0, dist_reg[224], 7'd0};
		4'd8: n_loc_oh_reg[31] = {7'd0, dist_reg[224], 8'd0};
		4'd9: n_loc_oh_reg[31] = {6'd0, dist_reg[224], 9'd0};
		4'd10: n_loc_oh_reg[31] = {5'd0, dist_reg[224], 10'd0};
		4'd11: n_loc_oh_reg[31] = {4'd0, dist_reg[224], 11'd0};
		4'd12: n_loc_oh_reg[31] = {3'd0, dist_reg[224], 12'd0};
		4'd13: n_loc_oh_reg[31] = {2'd0, dist_reg[224], 13'd0};
		4'd14: n_loc_oh_reg[31] = {1'd0, dist_reg[224], 14'd0};
		4'd15: n_loc_oh_reg[31] = {dist_reg[224], 15'd0};
	endcase
	case(loc_reg[32])
		4'd0: n_loc_oh_reg[32] = {15'd0, dist_reg[223]};
		4'd1: n_loc_oh_reg[32] = {14'd0, dist_reg[223], 1'd0};
		4'd2: n_loc_oh_reg[32] = {13'd0, dist_reg[223], 2'd0};
		4'd3: n_loc_oh_reg[32] = {12'd0, dist_reg[223], 3'd0};
		4'd4: n_loc_oh_reg[32] = {11'd0, dist_reg[223], 4'd0};
		4'd5: n_loc_oh_reg[32] = {10'd0, dist_reg[223], 5'd0};
		4'd6: n_loc_oh_reg[32] = {9'd0, dist_reg[223], 6'd0};
		4'd7: n_loc_oh_reg[32] = {8'd0, dist_reg[223], 7'd0};
		4'd8: n_loc_oh_reg[32] = {7'd0, dist_reg[223], 8'd0};
		4'd9: n_loc_oh_reg[32] = {6'd0, dist_reg[223], 9'd0};
		4'd10: n_loc_oh_reg[32] = {5'd0, dist_reg[223], 10'd0};
		4'd11: n_loc_oh_reg[32] = {4'd0, dist_reg[223], 11'd0};
		4'd12: n_loc_oh_reg[32] = {3'd0, dist_reg[223], 12'd0};
		4'd13: n_loc_oh_reg[32] = {2'd0, dist_reg[223], 13'd0};
		4'd14: n_loc_oh_reg[32] = {1'd0, dist_reg[223], 14'd0};
		4'd15: n_loc_oh_reg[32] = {dist_reg[223], 15'd0};
	endcase
	case(loc_reg[33])
		4'd0: n_loc_oh_reg[33] = {15'd0, dist_reg[222]};
		4'd1: n_loc_oh_reg[33] = {14'd0, dist_reg[222], 1'd0};
		4'd2: n_loc_oh_reg[33] = {13'd0, dist_reg[222], 2'd0};
		4'd3: n_loc_oh_reg[33] = {12'd0, dist_reg[222], 3'd0};
		4'd4: n_loc_oh_reg[33] = {11'd0, dist_reg[222], 4'd0};
		4'd5: n_loc_oh_reg[33] = {10'd0, dist_reg[222], 5'd0};
		4'd6: n_loc_oh_reg[33] = {9'd0, dist_reg[222], 6'd0};
		4'd7: n_loc_oh_reg[33] = {8'd0, dist_reg[222], 7'd0};
		4'd8: n_loc_oh_reg[33] = {7'd0, dist_reg[222], 8'd0};
		4'd9: n_loc_oh_reg[33] = {6'd0, dist_reg[222], 9'd0};
		4'd10: n_loc_oh_reg[33] = {5'd0, dist_reg[222], 10'd0};
		4'd11: n_loc_oh_reg[33] = {4'd0, dist_reg[222], 11'd0};
		4'd12: n_loc_oh_reg[33] = {3'd0, dist_reg[222], 12'd0};
		4'd13: n_loc_oh_reg[33] = {2'd0, dist_reg[222], 13'd0};
		4'd14: n_loc_oh_reg[33] = {1'd0, dist_reg[222], 14'd0};
		4'd15: n_loc_oh_reg[33] = {dist_reg[222], 15'd0};
	endcase
	case(loc_reg[34])
		4'd0: n_loc_oh_reg[34] = {15'd0, dist_reg[221]};
		4'd1: n_loc_oh_reg[34] = {14'd0, dist_reg[221], 1'd0};
		4'd2: n_loc_oh_reg[34] = {13'd0, dist_reg[221], 2'd0};
		4'd3: n_loc_oh_reg[34] = {12'd0, dist_reg[221], 3'd0};
		4'd4: n_loc_oh_reg[34] = {11'd0, dist_reg[221], 4'd0};
		4'd5: n_loc_oh_reg[34] = {10'd0, dist_reg[221], 5'd0};
		4'd6: n_loc_oh_reg[34] = {9'd0, dist_reg[221], 6'd0};
		4'd7: n_loc_oh_reg[34] = {8'd0, dist_reg[221], 7'd0};
		4'd8: n_loc_oh_reg[34] = {7'd0, dist_reg[221], 8'd0};
		4'd9: n_loc_oh_reg[34] = {6'd0, dist_reg[221], 9'd0};
		4'd10: n_loc_oh_reg[34] = {5'd0, dist_reg[221], 10'd0};
		4'd11: n_loc_oh_reg[34] = {4'd0, dist_reg[221], 11'd0};
		4'd12: n_loc_oh_reg[34] = {3'd0, dist_reg[221], 12'd0};
		4'd13: n_loc_oh_reg[34] = {2'd0, dist_reg[221], 13'd0};
		4'd14: n_loc_oh_reg[34] = {1'd0, dist_reg[221], 14'd0};
		4'd15: n_loc_oh_reg[34] = {dist_reg[221], 15'd0};
	endcase
	case(loc_reg[35])
		4'd0: n_loc_oh_reg[35] = {15'd0, dist_reg[220]};
		4'd1: n_loc_oh_reg[35] = {14'd0, dist_reg[220], 1'd0};
		4'd2: n_loc_oh_reg[35] = {13'd0, dist_reg[220], 2'd0};
		4'd3: n_loc_oh_reg[35] = {12'd0, dist_reg[220], 3'd0};
		4'd4: n_loc_oh_reg[35] = {11'd0, dist_reg[220], 4'd0};
		4'd5: n_loc_oh_reg[35] = {10'd0, dist_reg[220], 5'd0};
		4'd6: n_loc_oh_reg[35] = {9'd0, dist_reg[220], 6'd0};
		4'd7: n_loc_oh_reg[35] = {8'd0, dist_reg[220], 7'd0};
		4'd8: n_loc_oh_reg[35] = {7'd0, dist_reg[220], 8'd0};
		4'd9: n_loc_oh_reg[35] = {6'd0, dist_reg[220], 9'd0};
		4'd10: n_loc_oh_reg[35] = {5'd0, dist_reg[220], 10'd0};
		4'd11: n_loc_oh_reg[35] = {4'd0, dist_reg[220], 11'd0};
		4'd12: n_loc_oh_reg[35] = {3'd0, dist_reg[220], 12'd0};
		4'd13: n_loc_oh_reg[35] = {2'd0, dist_reg[220], 13'd0};
		4'd14: n_loc_oh_reg[35] = {1'd0, dist_reg[220], 14'd0};
		4'd15: n_loc_oh_reg[35] = {dist_reg[220], 15'd0};
	endcase
	case(loc_reg[36])
		4'd0: n_loc_oh_reg[36] = {15'd0, dist_reg[219]};
		4'd1: n_loc_oh_reg[36] = {14'd0, dist_reg[219], 1'd0};
		4'd2: n_loc_oh_reg[36] = {13'd0, dist_reg[219], 2'd0};
		4'd3: n_loc_oh_reg[36] = {12'd0, dist_reg[219], 3'd0};
		4'd4: n_loc_oh_reg[36] = {11'd0, dist_reg[219], 4'd0};
		4'd5: n_loc_oh_reg[36] = {10'd0, dist_reg[219], 5'd0};
		4'd6: n_loc_oh_reg[36] = {9'd0, dist_reg[219], 6'd0};
		4'd7: n_loc_oh_reg[36] = {8'd0, dist_reg[219], 7'd0};
		4'd8: n_loc_oh_reg[36] = {7'd0, dist_reg[219], 8'd0};
		4'd9: n_loc_oh_reg[36] = {6'd0, dist_reg[219], 9'd0};
		4'd10: n_loc_oh_reg[36] = {5'd0, dist_reg[219], 10'd0};
		4'd11: n_loc_oh_reg[36] = {4'd0, dist_reg[219], 11'd0};
		4'd12: n_loc_oh_reg[36] = {3'd0, dist_reg[219], 12'd0};
		4'd13: n_loc_oh_reg[36] = {2'd0, dist_reg[219], 13'd0};
		4'd14: n_loc_oh_reg[36] = {1'd0, dist_reg[219], 14'd0};
		4'd15: n_loc_oh_reg[36] = {dist_reg[219], 15'd0};
	endcase
	case(loc_reg[37])
		4'd0: n_loc_oh_reg[37] = {15'd0, dist_reg[218]};
		4'd1: n_loc_oh_reg[37] = {14'd0, dist_reg[218], 1'd0};
		4'd2: n_loc_oh_reg[37] = {13'd0, dist_reg[218], 2'd0};
		4'd3: n_loc_oh_reg[37] = {12'd0, dist_reg[218], 3'd0};
		4'd4: n_loc_oh_reg[37] = {11'd0, dist_reg[218], 4'd0};
		4'd5: n_loc_oh_reg[37] = {10'd0, dist_reg[218], 5'd0};
		4'd6: n_loc_oh_reg[37] = {9'd0, dist_reg[218], 6'd0};
		4'd7: n_loc_oh_reg[37] = {8'd0, dist_reg[218], 7'd0};
		4'd8: n_loc_oh_reg[37] = {7'd0, dist_reg[218], 8'd0};
		4'd9: n_loc_oh_reg[37] = {6'd0, dist_reg[218], 9'd0};
		4'd10: n_loc_oh_reg[37] = {5'd0, dist_reg[218], 10'd0};
		4'd11: n_loc_oh_reg[37] = {4'd0, dist_reg[218], 11'd0};
		4'd12: n_loc_oh_reg[37] = {3'd0, dist_reg[218], 12'd0};
		4'd13: n_loc_oh_reg[37] = {2'd0, dist_reg[218], 13'd0};
		4'd14: n_loc_oh_reg[37] = {1'd0, dist_reg[218], 14'd0};
		4'd15: n_loc_oh_reg[37] = {dist_reg[218], 15'd0};
	endcase
	case(loc_reg[38])
		4'd0: n_loc_oh_reg[38] = {15'd0, dist_reg[217]};
		4'd1: n_loc_oh_reg[38] = {14'd0, dist_reg[217], 1'd0};
		4'd2: n_loc_oh_reg[38] = {13'd0, dist_reg[217], 2'd0};
		4'd3: n_loc_oh_reg[38] = {12'd0, dist_reg[217], 3'd0};
		4'd4: n_loc_oh_reg[38] = {11'd0, dist_reg[217], 4'd0};
		4'd5: n_loc_oh_reg[38] = {10'd0, dist_reg[217], 5'd0};
		4'd6: n_loc_oh_reg[38] = {9'd0, dist_reg[217], 6'd0};
		4'd7: n_loc_oh_reg[38] = {8'd0, dist_reg[217], 7'd0};
		4'd8: n_loc_oh_reg[38] = {7'd0, dist_reg[217], 8'd0};
		4'd9: n_loc_oh_reg[38] = {6'd0, dist_reg[217], 9'd0};
		4'd10: n_loc_oh_reg[38] = {5'd0, dist_reg[217], 10'd0};
		4'd11: n_loc_oh_reg[38] = {4'd0, dist_reg[217], 11'd0};
		4'd12: n_loc_oh_reg[38] = {3'd0, dist_reg[217], 12'd0};
		4'd13: n_loc_oh_reg[38] = {2'd0, dist_reg[217], 13'd0};
		4'd14: n_loc_oh_reg[38] = {1'd0, dist_reg[217], 14'd0};
		4'd15: n_loc_oh_reg[38] = {dist_reg[217], 15'd0};
	endcase
	case(loc_reg[39])
		4'd0: n_loc_oh_reg[39] = {15'd0, dist_reg[216]};
		4'd1: n_loc_oh_reg[39] = {14'd0, dist_reg[216], 1'd0};
		4'd2: n_loc_oh_reg[39] = {13'd0, dist_reg[216], 2'd0};
		4'd3: n_loc_oh_reg[39] = {12'd0, dist_reg[216], 3'd0};
		4'd4: n_loc_oh_reg[39] = {11'd0, dist_reg[216], 4'd0};
		4'd5: n_loc_oh_reg[39] = {10'd0, dist_reg[216], 5'd0};
		4'd6: n_loc_oh_reg[39] = {9'd0, dist_reg[216], 6'd0};
		4'd7: n_loc_oh_reg[39] = {8'd0, dist_reg[216], 7'd0};
		4'd8: n_loc_oh_reg[39] = {7'd0, dist_reg[216], 8'd0};
		4'd9: n_loc_oh_reg[39] = {6'd0, dist_reg[216], 9'd0};
		4'd10: n_loc_oh_reg[39] = {5'd0, dist_reg[216], 10'd0};
		4'd11: n_loc_oh_reg[39] = {4'd0, dist_reg[216], 11'd0};
		4'd12: n_loc_oh_reg[39] = {3'd0, dist_reg[216], 12'd0};
		4'd13: n_loc_oh_reg[39] = {2'd0, dist_reg[216], 13'd0};
		4'd14: n_loc_oh_reg[39] = {1'd0, dist_reg[216], 14'd0};
		4'd15: n_loc_oh_reg[39] = {dist_reg[216], 15'd0};
	endcase
	case(loc_reg[40])
		4'd0: n_loc_oh_reg[40] = {15'd0, dist_reg[215]};
		4'd1: n_loc_oh_reg[40] = {14'd0, dist_reg[215], 1'd0};
		4'd2: n_loc_oh_reg[40] = {13'd0, dist_reg[215], 2'd0};
		4'd3: n_loc_oh_reg[40] = {12'd0, dist_reg[215], 3'd0};
		4'd4: n_loc_oh_reg[40] = {11'd0, dist_reg[215], 4'd0};
		4'd5: n_loc_oh_reg[40] = {10'd0, dist_reg[215], 5'd0};
		4'd6: n_loc_oh_reg[40] = {9'd0, dist_reg[215], 6'd0};
		4'd7: n_loc_oh_reg[40] = {8'd0, dist_reg[215], 7'd0};
		4'd8: n_loc_oh_reg[40] = {7'd0, dist_reg[215], 8'd0};
		4'd9: n_loc_oh_reg[40] = {6'd0, dist_reg[215], 9'd0};
		4'd10: n_loc_oh_reg[40] = {5'd0, dist_reg[215], 10'd0};
		4'd11: n_loc_oh_reg[40] = {4'd0, dist_reg[215], 11'd0};
		4'd12: n_loc_oh_reg[40] = {3'd0, dist_reg[215], 12'd0};
		4'd13: n_loc_oh_reg[40] = {2'd0, dist_reg[215], 13'd0};
		4'd14: n_loc_oh_reg[40] = {1'd0, dist_reg[215], 14'd0};
		4'd15: n_loc_oh_reg[40] = {dist_reg[215], 15'd0};
	endcase
	case(loc_reg[41])
		4'd0: n_loc_oh_reg[41] = {15'd0, dist_reg[214]};
		4'd1: n_loc_oh_reg[41] = {14'd0, dist_reg[214], 1'd0};
		4'd2: n_loc_oh_reg[41] = {13'd0, dist_reg[214], 2'd0};
		4'd3: n_loc_oh_reg[41] = {12'd0, dist_reg[214], 3'd0};
		4'd4: n_loc_oh_reg[41] = {11'd0, dist_reg[214], 4'd0};
		4'd5: n_loc_oh_reg[41] = {10'd0, dist_reg[214], 5'd0};
		4'd6: n_loc_oh_reg[41] = {9'd0, dist_reg[214], 6'd0};
		4'd7: n_loc_oh_reg[41] = {8'd0, dist_reg[214], 7'd0};
		4'd8: n_loc_oh_reg[41] = {7'd0, dist_reg[214], 8'd0};
		4'd9: n_loc_oh_reg[41] = {6'd0, dist_reg[214], 9'd0};
		4'd10: n_loc_oh_reg[41] = {5'd0, dist_reg[214], 10'd0};
		4'd11: n_loc_oh_reg[41] = {4'd0, dist_reg[214], 11'd0};
		4'd12: n_loc_oh_reg[41] = {3'd0, dist_reg[214], 12'd0};
		4'd13: n_loc_oh_reg[41] = {2'd0, dist_reg[214], 13'd0};
		4'd14: n_loc_oh_reg[41] = {1'd0, dist_reg[214], 14'd0};
		4'd15: n_loc_oh_reg[41] = {dist_reg[214], 15'd0};
	endcase
	case(loc_reg[42])
		4'd0: n_loc_oh_reg[42] = {15'd0, dist_reg[213]};
		4'd1: n_loc_oh_reg[42] = {14'd0, dist_reg[213], 1'd0};
		4'd2: n_loc_oh_reg[42] = {13'd0, dist_reg[213], 2'd0};
		4'd3: n_loc_oh_reg[42] = {12'd0, dist_reg[213], 3'd0};
		4'd4: n_loc_oh_reg[42] = {11'd0, dist_reg[213], 4'd0};
		4'd5: n_loc_oh_reg[42] = {10'd0, dist_reg[213], 5'd0};
		4'd6: n_loc_oh_reg[42] = {9'd0, dist_reg[213], 6'd0};
		4'd7: n_loc_oh_reg[42] = {8'd0, dist_reg[213], 7'd0};
		4'd8: n_loc_oh_reg[42] = {7'd0, dist_reg[213], 8'd0};
		4'd9: n_loc_oh_reg[42] = {6'd0, dist_reg[213], 9'd0};
		4'd10: n_loc_oh_reg[42] = {5'd0, dist_reg[213], 10'd0};
		4'd11: n_loc_oh_reg[42] = {4'd0, dist_reg[213], 11'd0};
		4'd12: n_loc_oh_reg[42] = {3'd0, dist_reg[213], 12'd0};
		4'd13: n_loc_oh_reg[42] = {2'd0, dist_reg[213], 13'd0};
		4'd14: n_loc_oh_reg[42] = {1'd0, dist_reg[213], 14'd0};
		4'd15: n_loc_oh_reg[42] = {dist_reg[213], 15'd0};
	endcase
	case(loc_reg[43])
		4'd0: n_loc_oh_reg[43] = {15'd0, dist_reg[212]};
		4'd1: n_loc_oh_reg[43] = {14'd0, dist_reg[212], 1'd0};
		4'd2: n_loc_oh_reg[43] = {13'd0, dist_reg[212], 2'd0};
		4'd3: n_loc_oh_reg[43] = {12'd0, dist_reg[212], 3'd0};
		4'd4: n_loc_oh_reg[43] = {11'd0, dist_reg[212], 4'd0};
		4'd5: n_loc_oh_reg[43] = {10'd0, dist_reg[212], 5'd0};
		4'd6: n_loc_oh_reg[43] = {9'd0, dist_reg[212], 6'd0};
		4'd7: n_loc_oh_reg[43] = {8'd0, dist_reg[212], 7'd0};
		4'd8: n_loc_oh_reg[43] = {7'd0, dist_reg[212], 8'd0};
		4'd9: n_loc_oh_reg[43] = {6'd0, dist_reg[212], 9'd0};
		4'd10: n_loc_oh_reg[43] = {5'd0, dist_reg[212], 10'd0};
		4'd11: n_loc_oh_reg[43] = {4'd0, dist_reg[212], 11'd0};
		4'd12: n_loc_oh_reg[43] = {3'd0, dist_reg[212], 12'd0};
		4'd13: n_loc_oh_reg[43] = {2'd0, dist_reg[212], 13'd0};
		4'd14: n_loc_oh_reg[43] = {1'd0, dist_reg[212], 14'd0};
		4'd15: n_loc_oh_reg[43] = {dist_reg[212], 15'd0};
	endcase
	case(loc_reg[44])
		4'd0: n_loc_oh_reg[44] = {15'd0, dist_reg[211]};
		4'd1: n_loc_oh_reg[44] = {14'd0, dist_reg[211], 1'd0};
		4'd2: n_loc_oh_reg[44] = {13'd0, dist_reg[211], 2'd0};
		4'd3: n_loc_oh_reg[44] = {12'd0, dist_reg[211], 3'd0};
		4'd4: n_loc_oh_reg[44] = {11'd0, dist_reg[211], 4'd0};
		4'd5: n_loc_oh_reg[44] = {10'd0, dist_reg[211], 5'd0};
		4'd6: n_loc_oh_reg[44] = {9'd0, dist_reg[211], 6'd0};
		4'd7: n_loc_oh_reg[44] = {8'd0, dist_reg[211], 7'd0};
		4'd8: n_loc_oh_reg[44] = {7'd0, dist_reg[211], 8'd0};
		4'd9: n_loc_oh_reg[44] = {6'd0, dist_reg[211], 9'd0};
		4'd10: n_loc_oh_reg[44] = {5'd0, dist_reg[211], 10'd0};
		4'd11: n_loc_oh_reg[44] = {4'd0, dist_reg[211], 11'd0};
		4'd12: n_loc_oh_reg[44] = {3'd0, dist_reg[211], 12'd0};
		4'd13: n_loc_oh_reg[44] = {2'd0, dist_reg[211], 13'd0};
		4'd14: n_loc_oh_reg[44] = {1'd0, dist_reg[211], 14'd0};
		4'd15: n_loc_oh_reg[44] = {dist_reg[211], 15'd0};
	endcase
	case(loc_reg[45])
		4'd0: n_loc_oh_reg[45] = {15'd0, dist_reg[210]};
		4'd1: n_loc_oh_reg[45] = {14'd0, dist_reg[210], 1'd0};
		4'd2: n_loc_oh_reg[45] = {13'd0, dist_reg[210], 2'd0};
		4'd3: n_loc_oh_reg[45] = {12'd0, dist_reg[210], 3'd0};
		4'd4: n_loc_oh_reg[45] = {11'd0, dist_reg[210], 4'd0};
		4'd5: n_loc_oh_reg[45] = {10'd0, dist_reg[210], 5'd0};
		4'd6: n_loc_oh_reg[45] = {9'd0, dist_reg[210], 6'd0};
		4'd7: n_loc_oh_reg[45] = {8'd0, dist_reg[210], 7'd0};
		4'd8: n_loc_oh_reg[45] = {7'd0, dist_reg[210], 8'd0};
		4'd9: n_loc_oh_reg[45] = {6'd0, dist_reg[210], 9'd0};
		4'd10: n_loc_oh_reg[45] = {5'd0, dist_reg[210], 10'd0};
		4'd11: n_loc_oh_reg[45] = {4'd0, dist_reg[210], 11'd0};
		4'd12: n_loc_oh_reg[45] = {3'd0, dist_reg[210], 12'd0};
		4'd13: n_loc_oh_reg[45] = {2'd0, dist_reg[210], 13'd0};
		4'd14: n_loc_oh_reg[45] = {1'd0, dist_reg[210], 14'd0};
		4'd15: n_loc_oh_reg[45] = {dist_reg[210], 15'd0};
	endcase
	case(loc_reg[46])
		4'd0: n_loc_oh_reg[46] = {15'd0, dist_reg[209]};
		4'd1: n_loc_oh_reg[46] = {14'd0, dist_reg[209], 1'd0};
		4'd2: n_loc_oh_reg[46] = {13'd0, dist_reg[209], 2'd0};
		4'd3: n_loc_oh_reg[46] = {12'd0, dist_reg[209], 3'd0};
		4'd4: n_loc_oh_reg[46] = {11'd0, dist_reg[209], 4'd0};
		4'd5: n_loc_oh_reg[46] = {10'd0, dist_reg[209], 5'd0};
		4'd6: n_loc_oh_reg[46] = {9'd0, dist_reg[209], 6'd0};
		4'd7: n_loc_oh_reg[46] = {8'd0, dist_reg[209], 7'd0};
		4'd8: n_loc_oh_reg[46] = {7'd0, dist_reg[209], 8'd0};
		4'd9: n_loc_oh_reg[46] = {6'd0, dist_reg[209], 9'd0};
		4'd10: n_loc_oh_reg[46] = {5'd0, dist_reg[209], 10'd0};
		4'd11: n_loc_oh_reg[46] = {4'd0, dist_reg[209], 11'd0};
		4'd12: n_loc_oh_reg[46] = {3'd0, dist_reg[209], 12'd0};
		4'd13: n_loc_oh_reg[46] = {2'd0, dist_reg[209], 13'd0};
		4'd14: n_loc_oh_reg[46] = {1'd0, dist_reg[209], 14'd0};
		4'd15: n_loc_oh_reg[46] = {dist_reg[209], 15'd0};
	endcase
	case(loc_reg[47])
		4'd0: n_loc_oh_reg[47] = {15'd0, dist_reg[208]};
		4'd1: n_loc_oh_reg[47] = {14'd0, dist_reg[208], 1'd0};
		4'd2: n_loc_oh_reg[47] = {13'd0, dist_reg[208], 2'd0};
		4'd3: n_loc_oh_reg[47] = {12'd0, dist_reg[208], 3'd0};
		4'd4: n_loc_oh_reg[47] = {11'd0, dist_reg[208], 4'd0};
		4'd5: n_loc_oh_reg[47] = {10'd0, dist_reg[208], 5'd0};
		4'd6: n_loc_oh_reg[47] = {9'd0, dist_reg[208], 6'd0};
		4'd7: n_loc_oh_reg[47] = {8'd0, dist_reg[208], 7'd0};
		4'd8: n_loc_oh_reg[47] = {7'd0, dist_reg[208], 8'd0};
		4'd9: n_loc_oh_reg[47] = {6'd0, dist_reg[208], 9'd0};
		4'd10: n_loc_oh_reg[47] = {5'd0, dist_reg[208], 10'd0};
		4'd11: n_loc_oh_reg[47] = {4'd0, dist_reg[208], 11'd0};
		4'd12: n_loc_oh_reg[47] = {3'd0, dist_reg[208], 12'd0};
		4'd13: n_loc_oh_reg[47] = {2'd0, dist_reg[208], 13'd0};
		4'd14: n_loc_oh_reg[47] = {1'd0, dist_reg[208], 14'd0};
		4'd15: n_loc_oh_reg[47] = {dist_reg[208], 15'd0};
	endcase
	case(loc_reg[48])
		4'd0: n_loc_oh_reg[48] = {15'd0, dist_reg[207]};
		4'd1: n_loc_oh_reg[48] = {14'd0, dist_reg[207], 1'd0};
		4'd2: n_loc_oh_reg[48] = {13'd0, dist_reg[207], 2'd0};
		4'd3: n_loc_oh_reg[48] = {12'd0, dist_reg[207], 3'd0};
		4'd4: n_loc_oh_reg[48] = {11'd0, dist_reg[207], 4'd0};
		4'd5: n_loc_oh_reg[48] = {10'd0, dist_reg[207], 5'd0};
		4'd6: n_loc_oh_reg[48] = {9'd0, dist_reg[207], 6'd0};
		4'd7: n_loc_oh_reg[48] = {8'd0, dist_reg[207], 7'd0};
		4'd8: n_loc_oh_reg[48] = {7'd0, dist_reg[207], 8'd0};
		4'd9: n_loc_oh_reg[48] = {6'd0, dist_reg[207], 9'd0};
		4'd10: n_loc_oh_reg[48] = {5'd0, dist_reg[207], 10'd0};
		4'd11: n_loc_oh_reg[48] = {4'd0, dist_reg[207], 11'd0};
		4'd12: n_loc_oh_reg[48] = {3'd0, dist_reg[207], 12'd0};
		4'd13: n_loc_oh_reg[48] = {2'd0, dist_reg[207], 13'd0};
		4'd14: n_loc_oh_reg[48] = {1'd0, dist_reg[207], 14'd0};
		4'd15: n_loc_oh_reg[48] = {dist_reg[207], 15'd0};
	endcase
	case(loc_reg[49])
		4'd0: n_loc_oh_reg[49] = {15'd0, dist_reg[206]};
		4'd1: n_loc_oh_reg[49] = {14'd0, dist_reg[206], 1'd0};
		4'd2: n_loc_oh_reg[49] = {13'd0, dist_reg[206], 2'd0};
		4'd3: n_loc_oh_reg[49] = {12'd0, dist_reg[206], 3'd0};
		4'd4: n_loc_oh_reg[49] = {11'd0, dist_reg[206], 4'd0};
		4'd5: n_loc_oh_reg[49] = {10'd0, dist_reg[206], 5'd0};
		4'd6: n_loc_oh_reg[49] = {9'd0, dist_reg[206], 6'd0};
		4'd7: n_loc_oh_reg[49] = {8'd0, dist_reg[206], 7'd0};
		4'd8: n_loc_oh_reg[49] = {7'd0, dist_reg[206], 8'd0};
		4'd9: n_loc_oh_reg[49] = {6'd0, dist_reg[206], 9'd0};
		4'd10: n_loc_oh_reg[49] = {5'd0, dist_reg[206], 10'd0};
		4'd11: n_loc_oh_reg[49] = {4'd0, dist_reg[206], 11'd0};
		4'd12: n_loc_oh_reg[49] = {3'd0, dist_reg[206], 12'd0};
		4'd13: n_loc_oh_reg[49] = {2'd0, dist_reg[206], 13'd0};
		4'd14: n_loc_oh_reg[49] = {1'd0, dist_reg[206], 14'd0};
		4'd15: n_loc_oh_reg[49] = {dist_reg[206], 15'd0};
	endcase
	case(loc_reg[50])
		4'd0: n_loc_oh_reg[50] = {15'd0, dist_reg[205]};
		4'd1: n_loc_oh_reg[50] = {14'd0, dist_reg[205], 1'd0};
		4'd2: n_loc_oh_reg[50] = {13'd0, dist_reg[205], 2'd0};
		4'd3: n_loc_oh_reg[50] = {12'd0, dist_reg[205], 3'd0};
		4'd4: n_loc_oh_reg[50] = {11'd0, dist_reg[205], 4'd0};
		4'd5: n_loc_oh_reg[50] = {10'd0, dist_reg[205], 5'd0};
		4'd6: n_loc_oh_reg[50] = {9'd0, dist_reg[205], 6'd0};
		4'd7: n_loc_oh_reg[50] = {8'd0, dist_reg[205], 7'd0};
		4'd8: n_loc_oh_reg[50] = {7'd0, dist_reg[205], 8'd0};
		4'd9: n_loc_oh_reg[50] = {6'd0, dist_reg[205], 9'd0};
		4'd10: n_loc_oh_reg[50] = {5'd0, dist_reg[205], 10'd0};
		4'd11: n_loc_oh_reg[50] = {4'd0, dist_reg[205], 11'd0};
		4'd12: n_loc_oh_reg[50] = {3'd0, dist_reg[205], 12'd0};
		4'd13: n_loc_oh_reg[50] = {2'd0, dist_reg[205], 13'd0};
		4'd14: n_loc_oh_reg[50] = {1'd0, dist_reg[205], 14'd0};
		4'd15: n_loc_oh_reg[50] = {dist_reg[205], 15'd0};
	endcase
	case(loc_reg[51])
		4'd0: n_loc_oh_reg[51] = {15'd0, dist_reg[204]};
		4'd1: n_loc_oh_reg[51] = {14'd0, dist_reg[204], 1'd0};
		4'd2: n_loc_oh_reg[51] = {13'd0, dist_reg[204], 2'd0};
		4'd3: n_loc_oh_reg[51] = {12'd0, dist_reg[204], 3'd0};
		4'd4: n_loc_oh_reg[51] = {11'd0, dist_reg[204], 4'd0};
		4'd5: n_loc_oh_reg[51] = {10'd0, dist_reg[204], 5'd0};
		4'd6: n_loc_oh_reg[51] = {9'd0, dist_reg[204], 6'd0};
		4'd7: n_loc_oh_reg[51] = {8'd0, dist_reg[204], 7'd0};
		4'd8: n_loc_oh_reg[51] = {7'd0, dist_reg[204], 8'd0};
		4'd9: n_loc_oh_reg[51] = {6'd0, dist_reg[204], 9'd0};
		4'd10: n_loc_oh_reg[51] = {5'd0, dist_reg[204], 10'd0};
		4'd11: n_loc_oh_reg[51] = {4'd0, dist_reg[204], 11'd0};
		4'd12: n_loc_oh_reg[51] = {3'd0, dist_reg[204], 12'd0};
		4'd13: n_loc_oh_reg[51] = {2'd0, dist_reg[204], 13'd0};
		4'd14: n_loc_oh_reg[51] = {1'd0, dist_reg[204], 14'd0};
		4'd15: n_loc_oh_reg[51] = {dist_reg[204], 15'd0};
	endcase
	case(loc_reg[52])
		4'd0: n_loc_oh_reg[52] = {15'd0, dist_reg[203]};
		4'd1: n_loc_oh_reg[52] = {14'd0, dist_reg[203], 1'd0};
		4'd2: n_loc_oh_reg[52] = {13'd0, dist_reg[203], 2'd0};
		4'd3: n_loc_oh_reg[52] = {12'd0, dist_reg[203], 3'd0};
		4'd4: n_loc_oh_reg[52] = {11'd0, dist_reg[203], 4'd0};
		4'd5: n_loc_oh_reg[52] = {10'd0, dist_reg[203], 5'd0};
		4'd6: n_loc_oh_reg[52] = {9'd0, dist_reg[203], 6'd0};
		4'd7: n_loc_oh_reg[52] = {8'd0, dist_reg[203], 7'd0};
		4'd8: n_loc_oh_reg[52] = {7'd0, dist_reg[203], 8'd0};
		4'd9: n_loc_oh_reg[52] = {6'd0, dist_reg[203], 9'd0};
		4'd10: n_loc_oh_reg[52] = {5'd0, dist_reg[203], 10'd0};
		4'd11: n_loc_oh_reg[52] = {4'd0, dist_reg[203], 11'd0};
		4'd12: n_loc_oh_reg[52] = {3'd0, dist_reg[203], 12'd0};
		4'd13: n_loc_oh_reg[52] = {2'd0, dist_reg[203], 13'd0};
		4'd14: n_loc_oh_reg[52] = {1'd0, dist_reg[203], 14'd0};
		4'd15: n_loc_oh_reg[52] = {dist_reg[203], 15'd0};
	endcase
	case(loc_reg[53])
		4'd0: n_loc_oh_reg[53] = {15'd0, dist_reg[202]};
		4'd1: n_loc_oh_reg[53] = {14'd0, dist_reg[202], 1'd0};
		4'd2: n_loc_oh_reg[53] = {13'd0, dist_reg[202], 2'd0};
		4'd3: n_loc_oh_reg[53] = {12'd0, dist_reg[202], 3'd0};
		4'd4: n_loc_oh_reg[53] = {11'd0, dist_reg[202], 4'd0};
		4'd5: n_loc_oh_reg[53] = {10'd0, dist_reg[202], 5'd0};
		4'd6: n_loc_oh_reg[53] = {9'd0, dist_reg[202], 6'd0};
		4'd7: n_loc_oh_reg[53] = {8'd0, dist_reg[202], 7'd0};
		4'd8: n_loc_oh_reg[53] = {7'd0, dist_reg[202], 8'd0};
		4'd9: n_loc_oh_reg[53] = {6'd0, dist_reg[202], 9'd0};
		4'd10: n_loc_oh_reg[53] = {5'd0, dist_reg[202], 10'd0};
		4'd11: n_loc_oh_reg[53] = {4'd0, dist_reg[202], 11'd0};
		4'd12: n_loc_oh_reg[53] = {3'd0, dist_reg[202], 12'd0};
		4'd13: n_loc_oh_reg[53] = {2'd0, dist_reg[202], 13'd0};
		4'd14: n_loc_oh_reg[53] = {1'd0, dist_reg[202], 14'd0};
		4'd15: n_loc_oh_reg[53] = {dist_reg[202], 15'd0};
	endcase
	case(loc_reg[54])
		4'd0: n_loc_oh_reg[54] = {15'd0, dist_reg[201]};
		4'd1: n_loc_oh_reg[54] = {14'd0, dist_reg[201], 1'd0};
		4'd2: n_loc_oh_reg[54] = {13'd0, dist_reg[201], 2'd0};
		4'd3: n_loc_oh_reg[54] = {12'd0, dist_reg[201], 3'd0};
		4'd4: n_loc_oh_reg[54] = {11'd0, dist_reg[201], 4'd0};
		4'd5: n_loc_oh_reg[54] = {10'd0, dist_reg[201], 5'd0};
		4'd6: n_loc_oh_reg[54] = {9'd0, dist_reg[201], 6'd0};
		4'd7: n_loc_oh_reg[54] = {8'd0, dist_reg[201], 7'd0};
		4'd8: n_loc_oh_reg[54] = {7'd0, dist_reg[201], 8'd0};
		4'd9: n_loc_oh_reg[54] = {6'd0, dist_reg[201], 9'd0};
		4'd10: n_loc_oh_reg[54] = {5'd0, dist_reg[201], 10'd0};
		4'd11: n_loc_oh_reg[54] = {4'd0, dist_reg[201], 11'd0};
		4'd12: n_loc_oh_reg[54] = {3'd0, dist_reg[201], 12'd0};
		4'd13: n_loc_oh_reg[54] = {2'd0, dist_reg[201], 13'd0};
		4'd14: n_loc_oh_reg[54] = {1'd0, dist_reg[201], 14'd0};
		4'd15: n_loc_oh_reg[54] = {dist_reg[201], 15'd0};
	endcase
	case(loc_reg[55])
		4'd0: n_loc_oh_reg[55] = {15'd0, dist_reg[200]};
		4'd1: n_loc_oh_reg[55] = {14'd0, dist_reg[200], 1'd0};
		4'd2: n_loc_oh_reg[55] = {13'd0, dist_reg[200], 2'd0};
		4'd3: n_loc_oh_reg[55] = {12'd0, dist_reg[200], 3'd0};
		4'd4: n_loc_oh_reg[55] = {11'd0, dist_reg[200], 4'd0};
		4'd5: n_loc_oh_reg[55] = {10'd0, dist_reg[200], 5'd0};
		4'd6: n_loc_oh_reg[55] = {9'd0, dist_reg[200], 6'd0};
		4'd7: n_loc_oh_reg[55] = {8'd0, dist_reg[200], 7'd0};
		4'd8: n_loc_oh_reg[55] = {7'd0, dist_reg[200], 8'd0};
		4'd9: n_loc_oh_reg[55] = {6'd0, dist_reg[200], 9'd0};
		4'd10: n_loc_oh_reg[55] = {5'd0, dist_reg[200], 10'd0};
		4'd11: n_loc_oh_reg[55] = {4'd0, dist_reg[200], 11'd0};
		4'd12: n_loc_oh_reg[55] = {3'd0, dist_reg[200], 12'd0};
		4'd13: n_loc_oh_reg[55] = {2'd0, dist_reg[200], 13'd0};
		4'd14: n_loc_oh_reg[55] = {1'd0, dist_reg[200], 14'd0};
		4'd15: n_loc_oh_reg[55] = {dist_reg[200], 15'd0};
	endcase
	case(loc_reg[56])
		4'd0: n_loc_oh_reg[56] = {15'd0, dist_reg[199]};
		4'd1: n_loc_oh_reg[56] = {14'd0, dist_reg[199], 1'd0};
		4'd2: n_loc_oh_reg[56] = {13'd0, dist_reg[199], 2'd0};
		4'd3: n_loc_oh_reg[56] = {12'd0, dist_reg[199], 3'd0};
		4'd4: n_loc_oh_reg[56] = {11'd0, dist_reg[199], 4'd0};
		4'd5: n_loc_oh_reg[56] = {10'd0, dist_reg[199], 5'd0};
		4'd6: n_loc_oh_reg[56] = {9'd0, dist_reg[199], 6'd0};
		4'd7: n_loc_oh_reg[56] = {8'd0, dist_reg[199], 7'd0};
		4'd8: n_loc_oh_reg[56] = {7'd0, dist_reg[199], 8'd0};
		4'd9: n_loc_oh_reg[56] = {6'd0, dist_reg[199], 9'd0};
		4'd10: n_loc_oh_reg[56] = {5'd0, dist_reg[199], 10'd0};
		4'd11: n_loc_oh_reg[56] = {4'd0, dist_reg[199], 11'd0};
		4'd12: n_loc_oh_reg[56] = {3'd0, dist_reg[199], 12'd0};
		4'd13: n_loc_oh_reg[56] = {2'd0, dist_reg[199], 13'd0};
		4'd14: n_loc_oh_reg[56] = {1'd0, dist_reg[199], 14'd0};
		4'd15: n_loc_oh_reg[56] = {dist_reg[199], 15'd0};
	endcase
	case(loc_reg[57])
		4'd0: n_loc_oh_reg[57] = {15'd0, dist_reg[198]};
		4'd1: n_loc_oh_reg[57] = {14'd0, dist_reg[198], 1'd0};
		4'd2: n_loc_oh_reg[57] = {13'd0, dist_reg[198], 2'd0};
		4'd3: n_loc_oh_reg[57] = {12'd0, dist_reg[198], 3'd0};
		4'd4: n_loc_oh_reg[57] = {11'd0, dist_reg[198], 4'd0};
		4'd5: n_loc_oh_reg[57] = {10'd0, dist_reg[198], 5'd0};
		4'd6: n_loc_oh_reg[57] = {9'd0, dist_reg[198], 6'd0};
		4'd7: n_loc_oh_reg[57] = {8'd0, dist_reg[198], 7'd0};
		4'd8: n_loc_oh_reg[57] = {7'd0, dist_reg[198], 8'd0};
		4'd9: n_loc_oh_reg[57] = {6'd0, dist_reg[198], 9'd0};
		4'd10: n_loc_oh_reg[57] = {5'd0, dist_reg[198], 10'd0};
		4'd11: n_loc_oh_reg[57] = {4'd0, dist_reg[198], 11'd0};
		4'd12: n_loc_oh_reg[57] = {3'd0, dist_reg[198], 12'd0};
		4'd13: n_loc_oh_reg[57] = {2'd0, dist_reg[198], 13'd0};
		4'd14: n_loc_oh_reg[57] = {1'd0, dist_reg[198], 14'd0};
		4'd15: n_loc_oh_reg[57] = {dist_reg[198], 15'd0};
	endcase
	case(loc_reg[58])
		4'd0: n_loc_oh_reg[58] = {15'd0, dist_reg[197]};
		4'd1: n_loc_oh_reg[58] = {14'd0, dist_reg[197], 1'd0};
		4'd2: n_loc_oh_reg[58] = {13'd0, dist_reg[197], 2'd0};
		4'd3: n_loc_oh_reg[58] = {12'd0, dist_reg[197], 3'd0};
		4'd4: n_loc_oh_reg[58] = {11'd0, dist_reg[197], 4'd0};
		4'd5: n_loc_oh_reg[58] = {10'd0, dist_reg[197], 5'd0};
		4'd6: n_loc_oh_reg[58] = {9'd0, dist_reg[197], 6'd0};
		4'd7: n_loc_oh_reg[58] = {8'd0, dist_reg[197], 7'd0};
		4'd8: n_loc_oh_reg[58] = {7'd0, dist_reg[197], 8'd0};
		4'd9: n_loc_oh_reg[58] = {6'd0, dist_reg[197], 9'd0};
		4'd10: n_loc_oh_reg[58] = {5'd0, dist_reg[197], 10'd0};
		4'd11: n_loc_oh_reg[58] = {4'd0, dist_reg[197], 11'd0};
		4'd12: n_loc_oh_reg[58] = {3'd0, dist_reg[197], 12'd0};
		4'd13: n_loc_oh_reg[58] = {2'd0, dist_reg[197], 13'd0};
		4'd14: n_loc_oh_reg[58] = {1'd0, dist_reg[197], 14'd0};
		4'd15: n_loc_oh_reg[58] = {dist_reg[197], 15'd0};
	endcase
	case(loc_reg[59])
		4'd0: n_loc_oh_reg[59] = {15'd0, dist_reg[196]};
		4'd1: n_loc_oh_reg[59] = {14'd0, dist_reg[196], 1'd0};
		4'd2: n_loc_oh_reg[59] = {13'd0, dist_reg[196], 2'd0};
		4'd3: n_loc_oh_reg[59] = {12'd0, dist_reg[196], 3'd0};
		4'd4: n_loc_oh_reg[59] = {11'd0, dist_reg[196], 4'd0};
		4'd5: n_loc_oh_reg[59] = {10'd0, dist_reg[196], 5'd0};
		4'd6: n_loc_oh_reg[59] = {9'd0, dist_reg[196], 6'd0};
		4'd7: n_loc_oh_reg[59] = {8'd0, dist_reg[196], 7'd0};
		4'd8: n_loc_oh_reg[59] = {7'd0, dist_reg[196], 8'd0};
		4'd9: n_loc_oh_reg[59] = {6'd0, dist_reg[196], 9'd0};
		4'd10: n_loc_oh_reg[59] = {5'd0, dist_reg[196], 10'd0};
		4'd11: n_loc_oh_reg[59] = {4'd0, dist_reg[196], 11'd0};
		4'd12: n_loc_oh_reg[59] = {3'd0, dist_reg[196], 12'd0};
		4'd13: n_loc_oh_reg[59] = {2'd0, dist_reg[196], 13'd0};
		4'd14: n_loc_oh_reg[59] = {1'd0, dist_reg[196], 14'd0};
		4'd15: n_loc_oh_reg[59] = {dist_reg[196], 15'd0};
	endcase
	case(loc_reg[60])
		4'd0: n_loc_oh_reg[60] = {15'd0, dist_reg[195]};
		4'd1: n_loc_oh_reg[60] = {14'd0, dist_reg[195], 1'd0};
		4'd2: n_loc_oh_reg[60] = {13'd0, dist_reg[195], 2'd0};
		4'd3: n_loc_oh_reg[60] = {12'd0, dist_reg[195], 3'd0};
		4'd4: n_loc_oh_reg[60] = {11'd0, dist_reg[195], 4'd0};
		4'd5: n_loc_oh_reg[60] = {10'd0, dist_reg[195], 5'd0};
		4'd6: n_loc_oh_reg[60] = {9'd0, dist_reg[195], 6'd0};
		4'd7: n_loc_oh_reg[60] = {8'd0, dist_reg[195], 7'd0};
		4'd8: n_loc_oh_reg[60] = {7'd0, dist_reg[195], 8'd0};
		4'd9: n_loc_oh_reg[60] = {6'd0, dist_reg[195], 9'd0};
		4'd10: n_loc_oh_reg[60] = {5'd0, dist_reg[195], 10'd0};
		4'd11: n_loc_oh_reg[60] = {4'd0, dist_reg[195], 11'd0};
		4'd12: n_loc_oh_reg[60] = {3'd0, dist_reg[195], 12'd0};
		4'd13: n_loc_oh_reg[60] = {2'd0, dist_reg[195], 13'd0};
		4'd14: n_loc_oh_reg[60] = {1'd0, dist_reg[195], 14'd0};
		4'd15: n_loc_oh_reg[60] = {dist_reg[195], 15'd0};
	endcase
	case(loc_reg[61])
		4'd0: n_loc_oh_reg[61] = {15'd0, dist_reg[194]};
		4'd1: n_loc_oh_reg[61] = {14'd0, dist_reg[194], 1'd0};
		4'd2: n_loc_oh_reg[61] = {13'd0, dist_reg[194], 2'd0};
		4'd3: n_loc_oh_reg[61] = {12'd0, dist_reg[194], 3'd0};
		4'd4: n_loc_oh_reg[61] = {11'd0, dist_reg[194], 4'd0};
		4'd5: n_loc_oh_reg[61] = {10'd0, dist_reg[194], 5'd0};
		4'd6: n_loc_oh_reg[61] = {9'd0, dist_reg[194], 6'd0};
		4'd7: n_loc_oh_reg[61] = {8'd0, dist_reg[194], 7'd0};
		4'd8: n_loc_oh_reg[61] = {7'd0, dist_reg[194], 8'd0};
		4'd9: n_loc_oh_reg[61] = {6'd0, dist_reg[194], 9'd0};
		4'd10: n_loc_oh_reg[61] = {5'd0, dist_reg[194], 10'd0};
		4'd11: n_loc_oh_reg[61] = {4'd0, dist_reg[194], 11'd0};
		4'd12: n_loc_oh_reg[61] = {3'd0, dist_reg[194], 12'd0};
		4'd13: n_loc_oh_reg[61] = {2'd0, dist_reg[194], 13'd0};
		4'd14: n_loc_oh_reg[61] = {1'd0, dist_reg[194], 14'd0};
		4'd15: n_loc_oh_reg[61] = {dist_reg[194], 15'd0};
	endcase
	case(loc_reg[62])
		4'd0: n_loc_oh_reg[62] = {15'd0, dist_reg[193]};
		4'd1: n_loc_oh_reg[62] = {14'd0, dist_reg[193], 1'd0};
		4'd2: n_loc_oh_reg[62] = {13'd0, dist_reg[193], 2'd0};
		4'd3: n_loc_oh_reg[62] = {12'd0, dist_reg[193], 3'd0};
		4'd4: n_loc_oh_reg[62] = {11'd0, dist_reg[193], 4'd0};
		4'd5: n_loc_oh_reg[62] = {10'd0, dist_reg[193], 5'd0};
		4'd6: n_loc_oh_reg[62] = {9'd0, dist_reg[193], 6'd0};
		4'd7: n_loc_oh_reg[62] = {8'd0, dist_reg[193], 7'd0};
		4'd8: n_loc_oh_reg[62] = {7'd0, dist_reg[193], 8'd0};
		4'd9: n_loc_oh_reg[62] = {6'd0, dist_reg[193], 9'd0};
		4'd10: n_loc_oh_reg[62] = {5'd0, dist_reg[193], 10'd0};
		4'd11: n_loc_oh_reg[62] = {4'd0, dist_reg[193], 11'd0};
		4'd12: n_loc_oh_reg[62] = {3'd0, dist_reg[193], 12'd0};
		4'd13: n_loc_oh_reg[62] = {2'd0, dist_reg[193], 13'd0};
		4'd14: n_loc_oh_reg[62] = {1'd0, dist_reg[193], 14'd0};
		4'd15: n_loc_oh_reg[62] = {dist_reg[193], 15'd0};
	endcase
	case(loc_reg[63])
		4'd0: n_loc_oh_reg[63] = {15'd0, dist_reg[192]};
		4'd1: n_loc_oh_reg[63] = {14'd0, dist_reg[192], 1'd0};
		4'd2: n_loc_oh_reg[63] = {13'd0, dist_reg[192], 2'd0};
		4'd3: n_loc_oh_reg[63] = {12'd0, dist_reg[192], 3'd0};
		4'd4: n_loc_oh_reg[63] = {11'd0, dist_reg[192], 4'd0};
		4'd5: n_loc_oh_reg[63] = {10'd0, dist_reg[192], 5'd0};
		4'd6: n_loc_oh_reg[63] = {9'd0, dist_reg[192], 6'd0};
		4'd7: n_loc_oh_reg[63] = {8'd0, dist_reg[192], 7'd0};
		4'd8: n_loc_oh_reg[63] = {7'd0, dist_reg[192], 8'd0};
		4'd9: n_loc_oh_reg[63] = {6'd0, dist_reg[192], 9'd0};
		4'd10: n_loc_oh_reg[63] = {5'd0, dist_reg[192], 10'd0};
		4'd11: n_loc_oh_reg[63] = {4'd0, dist_reg[192], 11'd0};
		4'd12: n_loc_oh_reg[63] = {3'd0, dist_reg[192], 12'd0};
		4'd13: n_loc_oh_reg[63] = {2'd0, dist_reg[192], 13'd0};
		4'd14: n_loc_oh_reg[63] = {1'd0, dist_reg[192], 14'd0};
		4'd15: n_loc_oh_reg[63] = {dist_reg[192], 15'd0};
	endcase
	case(loc_reg[64])
		4'd0: n_loc_oh_reg[64] = {15'd0, dist_reg[191]};
		4'd1: n_loc_oh_reg[64] = {14'd0, dist_reg[191], 1'd0};
		4'd2: n_loc_oh_reg[64] = {13'd0, dist_reg[191], 2'd0};
		4'd3: n_loc_oh_reg[64] = {12'd0, dist_reg[191], 3'd0};
		4'd4: n_loc_oh_reg[64] = {11'd0, dist_reg[191], 4'd0};
		4'd5: n_loc_oh_reg[64] = {10'd0, dist_reg[191], 5'd0};
		4'd6: n_loc_oh_reg[64] = {9'd0, dist_reg[191], 6'd0};
		4'd7: n_loc_oh_reg[64] = {8'd0, dist_reg[191], 7'd0};
		4'd8: n_loc_oh_reg[64] = {7'd0, dist_reg[191], 8'd0};
		4'd9: n_loc_oh_reg[64] = {6'd0, dist_reg[191], 9'd0};
		4'd10: n_loc_oh_reg[64] = {5'd0, dist_reg[191], 10'd0};
		4'd11: n_loc_oh_reg[64] = {4'd0, dist_reg[191], 11'd0};
		4'd12: n_loc_oh_reg[64] = {3'd0, dist_reg[191], 12'd0};
		4'd13: n_loc_oh_reg[64] = {2'd0, dist_reg[191], 13'd0};
		4'd14: n_loc_oh_reg[64] = {1'd0, dist_reg[191], 14'd0};
		4'd15: n_loc_oh_reg[64] = {dist_reg[191], 15'd0};
	endcase
	case(loc_reg[65])
		4'd0: n_loc_oh_reg[65] = {15'd0, dist_reg[190]};
		4'd1: n_loc_oh_reg[65] = {14'd0, dist_reg[190], 1'd0};
		4'd2: n_loc_oh_reg[65] = {13'd0, dist_reg[190], 2'd0};
		4'd3: n_loc_oh_reg[65] = {12'd0, dist_reg[190], 3'd0};
		4'd4: n_loc_oh_reg[65] = {11'd0, dist_reg[190], 4'd0};
		4'd5: n_loc_oh_reg[65] = {10'd0, dist_reg[190], 5'd0};
		4'd6: n_loc_oh_reg[65] = {9'd0, dist_reg[190], 6'd0};
		4'd7: n_loc_oh_reg[65] = {8'd0, dist_reg[190], 7'd0};
		4'd8: n_loc_oh_reg[65] = {7'd0, dist_reg[190], 8'd0};
		4'd9: n_loc_oh_reg[65] = {6'd0, dist_reg[190], 9'd0};
		4'd10: n_loc_oh_reg[65] = {5'd0, dist_reg[190], 10'd0};
		4'd11: n_loc_oh_reg[65] = {4'd0, dist_reg[190], 11'd0};
		4'd12: n_loc_oh_reg[65] = {3'd0, dist_reg[190], 12'd0};
		4'd13: n_loc_oh_reg[65] = {2'd0, dist_reg[190], 13'd0};
		4'd14: n_loc_oh_reg[65] = {1'd0, dist_reg[190], 14'd0};
		4'd15: n_loc_oh_reg[65] = {dist_reg[190], 15'd0};
	endcase
	case(loc_reg[66])
		4'd0: n_loc_oh_reg[66] = {15'd0, dist_reg[189]};
		4'd1: n_loc_oh_reg[66] = {14'd0, dist_reg[189], 1'd0};
		4'd2: n_loc_oh_reg[66] = {13'd0, dist_reg[189], 2'd0};
		4'd3: n_loc_oh_reg[66] = {12'd0, dist_reg[189], 3'd0};
		4'd4: n_loc_oh_reg[66] = {11'd0, dist_reg[189], 4'd0};
		4'd5: n_loc_oh_reg[66] = {10'd0, dist_reg[189], 5'd0};
		4'd6: n_loc_oh_reg[66] = {9'd0, dist_reg[189], 6'd0};
		4'd7: n_loc_oh_reg[66] = {8'd0, dist_reg[189], 7'd0};
		4'd8: n_loc_oh_reg[66] = {7'd0, dist_reg[189], 8'd0};
		4'd9: n_loc_oh_reg[66] = {6'd0, dist_reg[189], 9'd0};
		4'd10: n_loc_oh_reg[66] = {5'd0, dist_reg[189], 10'd0};
		4'd11: n_loc_oh_reg[66] = {4'd0, dist_reg[189], 11'd0};
		4'd12: n_loc_oh_reg[66] = {3'd0, dist_reg[189], 12'd0};
		4'd13: n_loc_oh_reg[66] = {2'd0, dist_reg[189], 13'd0};
		4'd14: n_loc_oh_reg[66] = {1'd0, dist_reg[189], 14'd0};
		4'd15: n_loc_oh_reg[66] = {dist_reg[189], 15'd0};
	endcase
	case(loc_reg[67])
		4'd0: n_loc_oh_reg[67] = {15'd0, dist_reg[188]};
		4'd1: n_loc_oh_reg[67] = {14'd0, dist_reg[188], 1'd0};
		4'd2: n_loc_oh_reg[67] = {13'd0, dist_reg[188], 2'd0};
		4'd3: n_loc_oh_reg[67] = {12'd0, dist_reg[188], 3'd0};
		4'd4: n_loc_oh_reg[67] = {11'd0, dist_reg[188], 4'd0};
		4'd5: n_loc_oh_reg[67] = {10'd0, dist_reg[188], 5'd0};
		4'd6: n_loc_oh_reg[67] = {9'd0, dist_reg[188], 6'd0};
		4'd7: n_loc_oh_reg[67] = {8'd0, dist_reg[188], 7'd0};
		4'd8: n_loc_oh_reg[67] = {7'd0, dist_reg[188], 8'd0};
		4'd9: n_loc_oh_reg[67] = {6'd0, dist_reg[188], 9'd0};
		4'd10: n_loc_oh_reg[67] = {5'd0, dist_reg[188], 10'd0};
		4'd11: n_loc_oh_reg[67] = {4'd0, dist_reg[188], 11'd0};
		4'd12: n_loc_oh_reg[67] = {3'd0, dist_reg[188], 12'd0};
		4'd13: n_loc_oh_reg[67] = {2'd0, dist_reg[188], 13'd0};
		4'd14: n_loc_oh_reg[67] = {1'd0, dist_reg[188], 14'd0};
		4'd15: n_loc_oh_reg[67] = {dist_reg[188], 15'd0};
	endcase
	case(loc_reg[68])
		4'd0: n_loc_oh_reg[68] = {15'd0, dist_reg[187]};
		4'd1: n_loc_oh_reg[68] = {14'd0, dist_reg[187], 1'd0};
		4'd2: n_loc_oh_reg[68] = {13'd0, dist_reg[187], 2'd0};
		4'd3: n_loc_oh_reg[68] = {12'd0, dist_reg[187], 3'd0};
		4'd4: n_loc_oh_reg[68] = {11'd0, dist_reg[187], 4'd0};
		4'd5: n_loc_oh_reg[68] = {10'd0, dist_reg[187], 5'd0};
		4'd6: n_loc_oh_reg[68] = {9'd0, dist_reg[187], 6'd0};
		4'd7: n_loc_oh_reg[68] = {8'd0, dist_reg[187], 7'd0};
		4'd8: n_loc_oh_reg[68] = {7'd0, dist_reg[187], 8'd0};
		4'd9: n_loc_oh_reg[68] = {6'd0, dist_reg[187], 9'd0};
		4'd10: n_loc_oh_reg[68] = {5'd0, dist_reg[187], 10'd0};
		4'd11: n_loc_oh_reg[68] = {4'd0, dist_reg[187], 11'd0};
		4'd12: n_loc_oh_reg[68] = {3'd0, dist_reg[187], 12'd0};
		4'd13: n_loc_oh_reg[68] = {2'd0, dist_reg[187], 13'd0};
		4'd14: n_loc_oh_reg[68] = {1'd0, dist_reg[187], 14'd0};
		4'd15: n_loc_oh_reg[68] = {dist_reg[187], 15'd0};
	endcase
	case(loc_reg[69])
		4'd0: n_loc_oh_reg[69] = {15'd0, dist_reg[186]};
		4'd1: n_loc_oh_reg[69] = {14'd0, dist_reg[186], 1'd0};
		4'd2: n_loc_oh_reg[69] = {13'd0, dist_reg[186], 2'd0};
		4'd3: n_loc_oh_reg[69] = {12'd0, dist_reg[186], 3'd0};
		4'd4: n_loc_oh_reg[69] = {11'd0, dist_reg[186], 4'd0};
		4'd5: n_loc_oh_reg[69] = {10'd0, dist_reg[186], 5'd0};
		4'd6: n_loc_oh_reg[69] = {9'd0, dist_reg[186], 6'd0};
		4'd7: n_loc_oh_reg[69] = {8'd0, dist_reg[186], 7'd0};
		4'd8: n_loc_oh_reg[69] = {7'd0, dist_reg[186], 8'd0};
		4'd9: n_loc_oh_reg[69] = {6'd0, dist_reg[186], 9'd0};
		4'd10: n_loc_oh_reg[69] = {5'd0, dist_reg[186], 10'd0};
		4'd11: n_loc_oh_reg[69] = {4'd0, dist_reg[186], 11'd0};
		4'd12: n_loc_oh_reg[69] = {3'd0, dist_reg[186], 12'd0};
		4'd13: n_loc_oh_reg[69] = {2'd0, dist_reg[186], 13'd0};
		4'd14: n_loc_oh_reg[69] = {1'd0, dist_reg[186], 14'd0};
		4'd15: n_loc_oh_reg[69] = {dist_reg[186], 15'd0};
	endcase
	case(loc_reg[70])
		4'd0: n_loc_oh_reg[70] = {15'd0, dist_reg[185]};
		4'd1: n_loc_oh_reg[70] = {14'd0, dist_reg[185], 1'd0};
		4'd2: n_loc_oh_reg[70] = {13'd0, dist_reg[185], 2'd0};
		4'd3: n_loc_oh_reg[70] = {12'd0, dist_reg[185], 3'd0};
		4'd4: n_loc_oh_reg[70] = {11'd0, dist_reg[185], 4'd0};
		4'd5: n_loc_oh_reg[70] = {10'd0, dist_reg[185], 5'd0};
		4'd6: n_loc_oh_reg[70] = {9'd0, dist_reg[185], 6'd0};
		4'd7: n_loc_oh_reg[70] = {8'd0, dist_reg[185], 7'd0};
		4'd8: n_loc_oh_reg[70] = {7'd0, dist_reg[185], 8'd0};
		4'd9: n_loc_oh_reg[70] = {6'd0, dist_reg[185], 9'd0};
		4'd10: n_loc_oh_reg[70] = {5'd0, dist_reg[185], 10'd0};
		4'd11: n_loc_oh_reg[70] = {4'd0, dist_reg[185], 11'd0};
		4'd12: n_loc_oh_reg[70] = {3'd0, dist_reg[185], 12'd0};
		4'd13: n_loc_oh_reg[70] = {2'd0, dist_reg[185], 13'd0};
		4'd14: n_loc_oh_reg[70] = {1'd0, dist_reg[185], 14'd0};
		4'd15: n_loc_oh_reg[70] = {dist_reg[185], 15'd0};
	endcase
	case(loc_reg[71])
		4'd0: n_loc_oh_reg[71] = {15'd0, dist_reg[184]};
		4'd1: n_loc_oh_reg[71] = {14'd0, dist_reg[184], 1'd0};
		4'd2: n_loc_oh_reg[71] = {13'd0, dist_reg[184], 2'd0};
		4'd3: n_loc_oh_reg[71] = {12'd0, dist_reg[184], 3'd0};
		4'd4: n_loc_oh_reg[71] = {11'd0, dist_reg[184], 4'd0};
		4'd5: n_loc_oh_reg[71] = {10'd0, dist_reg[184], 5'd0};
		4'd6: n_loc_oh_reg[71] = {9'd0, dist_reg[184], 6'd0};
		4'd7: n_loc_oh_reg[71] = {8'd0, dist_reg[184], 7'd0};
		4'd8: n_loc_oh_reg[71] = {7'd0, dist_reg[184], 8'd0};
		4'd9: n_loc_oh_reg[71] = {6'd0, dist_reg[184], 9'd0};
		4'd10: n_loc_oh_reg[71] = {5'd0, dist_reg[184], 10'd0};
		4'd11: n_loc_oh_reg[71] = {4'd0, dist_reg[184], 11'd0};
		4'd12: n_loc_oh_reg[71] = {3'd0, dist_reg[184], 12'd0};
		4'd13: n_loc_oh_reg[71] = {2'd0, dist_reg[184], 13'd0};
		4'd14: n_loc_oh_reg[71] = {1'd0, dist_reg[184], 14'd0};
		4'd15: n_loc_oh_reg[71] = {dist_reg[184], 15'd0};
	endcase
	case(loc_reg[72])
		4'd0: n_loc_oh_reg[72] = {15'd0, dist_reg[183]};
		4'd1: n_loc_oh_reg[72] = {14'd0, dist_reg[183], 1'd0};
		4'd2: n_loc_oh_reg[72] = {13'd0, dist_reg[183], 2'd0};
		4'd3: n_loc_oh_reg[72] = {12'd0, dist_reg[183], 3'd0};
		4'd4: n_loc_oh_reg[72] = {11'd0, dist_reg[183], 4'd0};
		4'd5: n_loc_oh_reg[72] = {10'd0, dist_reg[183], 5'd0};
		4'd6: n_loc_oh_reg[72] = {9'd0, dist_reg[183], 6'd0};
		4'd7: n_loc_oh_reg[72] = {8'd0, dist_reg[183], 7'd0};
		4'd8: n_loc_oh_reg[72] = {7'd0, dist_reg[183], 8'd0};
		4'd9: n_loc_oh_reg[72] = {6'd0, dist_reg[183], 9'd0};
		4'd10: n_loc_oh_reg[72] = {5'd0, dist_reg[183], 10'd0};
		4'd11: n_loc_oh_reg[72] = {4'd0, dist_reg[183], 11'd0};
		4'd12: n_loc_oh_reg[72] = {3'd0, dist_reg[183], 12'd0};
		4'd13: n_loc_oh_reg[72] = {2'd0, dist_reg[183], 13'd0};
		4'd14: n_loc_oh_reg[72] = {1'd0, dist_reg[183], 14'd0};
		4'd15: n_loc_oh_reg[72] = {dist_reg[183], 15'd0};
	endcase
	case(loc_reg[73])
		4'd0: n_loc_oh_reg[73] = {15'd0, dist_reg[182]};
		4'd1: n_loc_oh_reg[73] = {14'd0, dist_reg[182], 1'd0};
		4'd2: n_loc_oh_reg[73] = {13'd0, dist_reg[182], 2'd0};
		4'd3: n_loc_oh_reg[73] = {12'd0, dist_reg[182], 3'd0};
		4'd4: n_loc_oh_reg[73] = {11'd0, dist_reg[182], 4'd0};
		4'd5: n_loc_oh_reg[73] = {10'd0, dist_reg[182], 5'd0};
		4'd6: n_loc_oh_reg[73] = {9'd0, dist_reg[182], 6'd0};
		4'd7: n_loc_oh_reg[73] = {8'd0, dist_reg[182], 7'd0};
		4'd8: n_loc_oh_reg[73] = {7'd0, dist_reg[182], 8'd0};
		4'd9: n_loc_oh_reg[73] = {6'd0, dist_reg[182], 9'd0};
		4'd10: n_loc_oh_reg[73] = {5'd0, dist_reg[182], 10'd0};
		4'd11: n_loc_oh_reg[73] = {4'd0, dist_reg[182], 11'd0};
		4'd12: n_loc_oh_reg[73] = {3'd0, dist_reg[182], 12'd0};
		4'd13: n_loc_oh_reg[73] = {2'd0, dist_reg[182], 13'd0};
		4'd14: n_loc_oh_reg[73] = {1'd0, dist_reg[182], 14'd0};
		4'd15: n_loc_oh_reg[73] = {dist_reg[182], 15'd0};
	endcase
	case(loc_reg[74])
		4'd0: n_loc_oh_reg[74] = {15'd0, dist_reg[181]};
		4'd1: n_loc_oh_reg[74] = {14'd0, dist_reg[181], 1'd0};
		4'd2: n_loc_oh_reg[74] = {13'd0, dist_reg[181], 2'd0};
		4'd3: n_loc_oh_reg[74] = {12'd0, dist_reg[181], 3'd0};
		4'd4: n_loc_oh_reg[74] = {11'd0, dist_reg[181], 4'd0};
		4'd5: n_loc_oh_reg[74] = {10'd0, dist_reg[181], 5'd0};
		4'd6: n_loc_oh_reg[74] = {9'd0, dist_reg[181], 6'd0};
		4'd7: n_loc_oh_reg[74] = {8'd0, dist_reg[181], 7'd0};
		4'd8: n_loc_oh_reg[74] = {7'd0, dist_reg[181], 8'd0};
		4'd9: n_loc_oh_reg[74] = {6'd0, dist_reg[181], 9'd0};
		4'd10: n_loc_oh_reg[74] = {5'd0, dist_reg[181], 10'd0};
		4'd11: n_loc_oh_reg[74] = {4'd0, dist_reg[181], 11'd0};
		4'd12: n_loc_oh_reg[74] = {3'd0, dist_reg[181], 12'd0};
		4'd13: n_loc_oh_reg[74] = {2'd0, dist_reg[181], 13'd0};
		4'd14: n_loc_oh_reg[74] = {1'd0, dist_reg[181], 14'd0};
		4'd15: n_loc_oh_reg[74] = {dist_reg[181], 15'd0};
	endcase
	case(loc_reg[75])
		4'd0: n_loc_oh_reg[75] = {15'd0, dist_reg[180]};
		4'd1: n_loc_oh_reg[75] = {14'd0, dist_reg[180], 1'd0};
		4'd2: n_loc_oh_reg[75] = {13'd0, dist_reg[180], 2'd0};
		4'd3: n_loc_oh_reg[75] = {12'd0, dist_reg[180], 3'd0};
		4'd4: n_loc_oh_reg[75] = {11'd0, dist_reg[180], 4'd0};
		4'd5: n_loc_oh_reg[75] = {10'd0, dist_reg[180], 5'd0};
		4'd6: n_loc_oh_reg[75] = {9'd0, dist_reg[180], 6'd0};
		4'd7: n_loc_oh_reg[75] = {8'd0, dist_reg[180], 7'd0};
		4'd8: n_loc_oh_reg[75] = {7'd0, dist_reg[180], 8'd0};
		4'd9: n_loc_oh_reg[75] = {6'd0, dist_reg[180], 9'd0};
		4'd10: n_loc_oh_reg[75] = {5'd0, dist_reg[180], 10'd0};
		4'd11: n_loc_oh_reg[75] = {4'd0, dist_reg[180], 11'd0};
		4'd12: n_loc_oh_reg[75] = {3'd0, dist_reg[180], 12'd0};
		4'd13: n_loc_oh_reg[75] = {2'd0, dist_reg[180], 13'd0};
		4'd14: n_loc_oh_reg[75] = {1'd0, dist_reg[180], 14'd0};
		4'd15: n_loc_oh_reg[75] = {dist_reg[180], 15'd0};
	endcase
	case(loc_reg[76])
		4'd0: n_loc_oh_reg[76] = {15'd0, dist_reg[179]};
		4'd1: n_loc_oh_reg[76] = {14'd0, dist_reg[179], 1'd0};
		4'd2: n_loc_oh_reg[76] = {13'd0, dist_reg[179], 2'd0};
		4'd3: n_loc_oh_reg[76] = {12'd0, dist_reg[179], 3'd0};
		4'd4: n_loc_oh_reg[76] = {11'd0, dist_reg[179], 4'd0};
		4'd5: n_loc_oh_reg[76] = {10'd0, dist_reg[179], 5'd0};
		4'd6: n_loc_oh_reg[76] = {9'd0, dist_reg[179], 6'd0};
		4'd7: n_loc_oh_reg[76] = {8'd0, dist_reg[179], 7'd0};
		4'd8: n_loc_oh_reg[76] = {7'd0, dist_reg[179], 8'd0};
		4'd9: n_loc_oh_reg[76] = {6'd0, dist_reg[179], 9'd0};
		4'd10: n_loc_oh_reg[76] = {5'd0, dist_reg[179], 10'd0};
		4'd11: n_loc_oh_reg[76] = {4'd0, dist_reg[179], 11'd0};
		4'd12: n_loc_oh_reg[76] = {3'd0, dist_reg[179], 12'd0};
		4'd13: n_loc_oh_reg[76] = {2'd0, dist_reg[179], 13'd0};
		4'd14: n_loc_oh_reg[76] = {1'd0, dist_reg[179], 14'd0};
		4'd15: n_loc_oh_reg[76] = {dist_reg[179], 15'd0};
	endcase
	case(loc_reg[77])
		4'd0: n_loc_oh_reg[77] = {15'd0, dist_reg[178]};
		4'd1: n_loc_oh_reg[77] = {14'd0, dist_reg[178], 1'd0};
		4'd2: n_loc_oh_reg[77] = {13'd0, dist_reg[178], 2'd0};
		4'd3: n_loc_oh_reg[77] = {12'd0, dist_reg[178], 3'd0};
		4'd4: n_loc_oh_reg[77] = {11'd0, dist_reg[178], 4'd0};
		4'd5: n_loc_oh_reg[77] = {10'd0, dist_reg[178], 5'd0};
		4'd6: n_loc_oh_reg[77] = {9'd0, dist_reg[178], 6'd0};
		4'd7: n_loc_oh_reg[77] = {8'd0, dist_reg[178], 7'd0};
		4'd8: n_loc_oh_reg[77] = {7'd0, dist_reg[178], 8'd0};
		4'd9: n_loc_oh_reg[77] = {6'd0, dist_reg[178], 9'd0};
		4'd10: n_loc_oh_reg[77] = {5'd0, dist_reg[178], 10'd0};
		4'd11: n_loc_oh_reg[77] = {4'd0, dist_reg[178], 11'd0};
		4'd12: n_loc_oh_reg[77] = {3'd0, dist_reg[178], 12'd0};
		4'd13: n_loc_oh_reg[77] = {2'd0, dist_reg[178], 13'd0};
		4'd14: n_loc_oh_reg[77] = {1'd0, dist_reg[178], 14'd0};
		4'd15: n_loc_oh_reg[77] = {dist_reg[178], 15'd0};
	endcase
	case(loc_reg[78])
		4'd0: n_loc_oh_reg[78] = {15'd0, dist_reg[177]};
		4'd1: n_loc_oh_reg[78] = {14'd0, dist_reg[177], 1'd0};
		4'd2: n_loc_oh_reg[78] = {13'd0, dist_reg[177], 2'd0};
		4'd3: n_loc_oh_reg[78] = {12'd0, dist_reg[177], 3'd0};
		4'd4: n_loc_oh_reg[78] = {11'd0, dist_reg[177], 4'd0};
		4'd5: n_loc_oh_reg[78] = {10'd0, dist_reg[177], 5'd0};
		4'd6: n_loc_oh_reg[78] = {9'd0, dist_reg[177], 6'd0};
		4'd7: n_loc_oh_reg[78] = {8'd0, dist_reg[177], 7'd0};
		4'd8: n_loc_oh_reg[78] = {7'd0, dist_reg[177], 8'd0};
		4'd9: n_loc_oh_reg[78] = {6'd0, dist_reg[177], 9'd0};
		4'd10: n_loc_oh_reg[78] = {5'd0, dist_reg[177], 10'd0};
		4'd11: n_loc_oh_reg[78] = {4'd0, dist_reg[177], 11'd0};
		4'd12: n_loc_oh_reg[78] = {3'd0, dist_reg[177], 12'd0};
		4'd13: n_loc_oh_reg[78] = {2'd0, dist_reg[177], 13'd0};
		4'd14: n_loc_oh_reg[78] = {1'd0, dist_reg[177], 14'd0};
		4'd15: n_loc_oh_reg[78] = {dist_reg[177], 15'd0};
	endcase
	case(loc_reg[79])
		4'd0: n_loc_oh_reg[79] = {15'd0, dist_reg[176]};
		4'd1: n_loc_oh_reg[79] = {14'd0, dist_reg[176], 1'd0};
		4'd2: n_loc_oh_reg[79] = {13'd0, dist_reg[176], 2'd0};
		4'd3: n_loc_oh_reg[79] = {12'd0, dist_reg[176], 3'd0};
		4'd4: n_loc_oh_reg[79] = {11'd0, dist_reg[176], 4'd0};
		4'd5: n_loc_oh_reg[79] = {10'd0, dist_reg[176], 5'd0};
		4'd6: n_loc_oh_reg[79] = {9'd0, dist_reg[176], 6'd0};
		4'd7: n_loc_oh_reg[79] = {8'd0, dist_reg[176], 7'd0};
		4'd8: n_loc_oh_reg[79] = {7'd0, dist_reg[176], 8'd0};
		4'd9: n_loc_oh_reg[79] = {6'd0, dist_reg[176], 9'd0};
		4'd10: n_loc_oh_reg[79] = {5'd0, dist_reg[176], 10'd0};
		4'd11: n_loc_oh_reg[79] = {4'd0, dist_reg[176], 11'd0};
		4'd12: n_loc_oh_reg[79] = {3'd0, dist_reg[176], 12'd0};
		4'd13: n_loc_oh_reg[79] = {2'd0, dist_reg[176], 13'd0};
		4'd14: n_loc_oh_reg[79] = {1'd0, dist_reg[176], 14'd0};
		4'd15: n_loc_oh_reg[79] = {dist_reg[176], 15'd0};
	endcase
	case(loc_reg[80])
		4'd0: n_loc_oh_reg[80] = {15'd0, dist_reg[175]};
		4'd1: n_loc_oh_reg[80] = {14'd0, dist_reg[175], 1'd0};
		4'd2: n_loc_oh_reg[80] = {13'd0, dist_reg[175], 2'd0};
		4'd3: n_loc_oh_reg[80] = {12'd0, dist_reg[175], 3'd0};
		4'd4: n_loc_oh_reg[80] = {11'd0, dist_reg[175], 4'd0};
		4'd5: n_loc_oh_reg[80] = {10'd0, dist_reg[175], 5'd0};
		4'd6: n_loc_oh_reg[80] = {9'd0, dist_reg[175], 6'd0};
		4'd7: n_loc_oh_reg[80] = {8'd0, dist_reg[175], 7'd0};
		4'd8: n_loc_oh_reg[80] = {7'd0, dist_reg[175], 8'd0};
		4'd9: n_loc_oh_reg[80] = {6'd0, dist_reg[175], 9'd0};
		4'd10: n_loc_oh_reg[80] = {5'd0, dist_reg[175], 10'd0};
		4'd11: n_loc_oh_reg[80] = {4'd0, dist_reg[175], 11'd0};
		4'd12: n_loc_oh_reg[80] = {3'd0, dist_reg[175], 12'd0};
		4'd13: n_loc_oh_reg[80] = {2'd0, dist_reg[175], 13'd0};
		4'd14: n_loc_oh_reg[80] = {1'd0, dist_reg[175], 14'd0};
		4'd15: n_loc_oh_reg[80] = {dist_reg[175], 15'd0};
	endcase
	case(loc_reg[81])
		4'd0: n_loc_oh_reg[81] = {15'd0, dist_reg[174]};
		4'd1: n_loc_oh_reg[81] = {14'd0, dist_reg[174], 1'd0};
		4'd2: n_loc_oh_reg[81] = {13'd0, dist_reg[174], 2'd0};
		4'd3: n_loc_oh_reg[81] = {12'd0, dist_reg[174], 3'd0};
		4'd4: n_loc_oh_reg[81] = {11'd0, dist_reg[174], 4'd0};
		4'd5: n_loc_oh_reg[81] = {10'd0, dist_reg[174], 5'd0};
		4'd6: n_loc_oh_reg[81] = {9'd0, dist_reg[174], 6'd0};
		4'd7: n_loc_oh_reg[81] = {8'd0, dist_reg[174], 7'd0};
		4'd8: n_loc_oh_reg[81] = {7'd0, dist_reg[174], 8'd0};
		4'd9: n_loc_oh_reg[81] = {6'd0, dist_reg[174], 9'd0};
		4'd10: n_loc_oh_reg[81] = {5'd0, dist_reg[174], 10'd0};
		4'd11: n_loc_oh_reg[81] = {4'd0, dist_reg[174], 11'd0};
		4'd12: n_loc_oh_reg[81] = {3'd0, dist_reg[174], 12'd0};
		4'd13: n_loc_oh_reg[81] = {2'd0, dist_reg[174], 13'd0};
		4'd14: n_loc_oh_reg[81] = {1'd0, dist_reg[174], 14'd0};
		4'd15: n_loc_oh_reg[81] = {dist_reg[174], 15'd0};
	endcase
	case(loc_reg[82])
		4'd0: n_loc_oh_reg[82] = {15'd0, dist_reg[173]};
		4'd1: n_loc_oh_reg[82] = {14'd0, dist_reg[173], 1'd0};
		4'd2: n_loc_oh_reg[82] = {13'd0, dist_reg[173], 2'd0};
		4'd3: n_loc_oh_reg[82] = {12'd0, dist_reg[173], 3'd0};
		4'd4: n_loc_oh_reg[82] = {11'd0, dist_reg[173], 4'd0};
		4'd5: n_loc_oh_reg[82] = {10'd0, dist_reg[173], 5'd0};
		4'd6: n_loc_oh_reg[82] = {9'd0, dist_reg[173], 6'd0};
		4'd7: n_loc_oh_reg[82] = {8'd0, dist_reg[173], 7'd0};
		4'd8: n_loc_oh_reg[82] = {7'd0, dist_reg[173], 8'd0};
		4'd9: n_loc_oh_reg[82] = {6'd0, dist_reg[173], 9'd0};
		4'd10: n_loc_oh_reg[82] = {5'd0, dist_reg[173], 10'd0};
		4'd11: n_loc_oh_reg[82] = {4'd0, dist_reg[173], 11'd0};
		4'd12: n_loc_oh_reg[82] = {3'd0, dist_reg[173], 12'd0};
		4'd13: n_loc_oh_reg[82] = {2'd0, dist_reg[173], 13'd0};
		4'd14: n_loc_oh_reg[82] = {1'd0, dist_reg[173], 14'd0};
		4'd15: n_loc_oh_reg[82] = {dist_reg[173], 15'd0};
	endcase
	case(loc_reg[83])
		4'd0: n_loc_oh_reg[83] = {15'd0, dist_reg[172]};
		4'd1: n_loc_oh_reg[83] = {14'd0, dist_reg[172], 1'd0};
		4'd2: n_loc_oh_reg[83] = {13'd0, dist_reg[172], 2'd0};
		4'd3: n_loc_oh_reg[83] = {12'd0, dist_reg[172], 3'd0};
		4'd4: n_loc_oh_reg[83] = {11'd0, dist_reg[172], 4'd0};
		4'd5: n_loc_oh_reg[83] = {10'd0, dist_reg[172], 5'd0};
		4'd6: n_loc_oh_reg[83] = {9'd0, dist_reg[172], 6'd0};
		4'd7: n_loc_oh_reg[83] = {8'd0, dist_reg[172], 7'd0};
		4'd8: n_loc_oh_reg[83] = {7'd0, dist_reg[172], 8'd0};
		4'd9: n_loc_oh_reg[83] = {6'd0, dist_reg[172], 9'd0};
		4'd10: n_loc_oh_reg[83] = {5'd0, dist_reg[172], 10'd0};
		4'd11: n_loc_oh_reg[83] = {4'd0, dist_reg[172], 11'd0};
		4'd12: n_loc_oh_reg[83] = {3'd0, dist_reg[172], 12'd0};
		4'd13: n_loc_oh_reg[83] = {2'd0, dist_reg[172], 13'd0};
		4'd14: n_loc_oh_reg[83] = {1'd0, dist_reg[172], 14'd0};
		4'd15: n_loc_oh_reg[83] = {dist_reg[172], 15'd0};
	endcase
	case(loc_reg[84])
		4'd0: n_loc_oh_reg[84] = {15'd0, dist_reg[171]};
		4'd1: n_loc_oh_reg[84] = {14'd0, dist_reg[171], 1'd0};
		4'd2: n_loc_oh_reg[84] = {13'd0, dist_reg[171], 2'd0};
		4'd3: n_loc_oh_reg[84] = {12'd0, dist_reg[171], 3'd0};
		4'd4: n_loc_oh_reg[84] = {11'd0, dist_reg[171], 4'd0};
		4'd5: n_loc_oh_reg[84] = {10'd0, dist_reg[171], 5'd0};
		4'd6: n_loc_oh_reg[84] = {9'd0, dist_reg[171], 6'd0};
		4'd7: n_loc_oh_reg[84] = {8'd0, dist_reg[171], 7'd0};
		4'd8: n_loc_oh_reg[84] = {7'd0, dist_reg[171], 8'd0};
		4'd9: n_loc_oh_reg[84] = {6'd0, dist_reg[171], 9'd0};
		4'd10: n_loc_oh_reg[84] = {5'd0, dist_reg[171], 10'd0};
		4'd11: n_loc_oh_reg[84] = {4'd0, dist_reg[171], 11'd0};
		4'd12: n_loc_oh_reg[84] = {3'd0, dist_reg[171], 12'd0};
		4'd13: n_loc_oh_reg[84] = {2'd0, dist_reg[171], 13'd0};
		4'd14: n_loc_oh_reg[84] = {1'd0, dist_reg[171], 14'd0};
		4'd15: n_loc_oh_reg[84] = {dist_reg[171], 15'd0};
	endcase
	case(loc_reg[85])
		4'd0: n_loc_oh_reg[85] = {15'd0, dist_reg[170]};
		4'd1: n_loc_oh_reg[85] = {14'd0, dist_reg[170], 1'd0};
		4'd2: n_loc_oh_reg[85] = {13'd0, dist_reg[170], 2'd0};
		4'd3: n_loc_oh_reg[85] = {12'd0, dist_reg[170], 3'd0};
		4'd4: n_loc_oh_reg[85] = {11'd0, dist_reg[170], 4'd0};
		4'd5: n_loc_oh_reg[85] = {10'd0, dist_reg[170], 5'd0};
		4'd6: n_loc_oh_reg[85] = {9'd0, dist_reg[170], 6'd0};
		4'd7: n_loc_oh_reg[85] = {8'd0, dist_reg[170], 7'd0};
		4'd8: n_loc_oh_reg[85] = {7'd0, dist_reg[170], 8'd0};
		4'd9: n_loc_oh_reg[85] = {6'd0, dist_reg[170], 9'd0};
		4'd10: n_loc_oh_reg[85] = {5'd0, dist_reg[170], 10'd0};
		4'd11: n_loc_oh_reg[85] = {4'd0, dist_reg[170], 11'd0};
		4'd12: n_loc_oh_reg[85] = {3'd0, dist_reg[170], 12'd0};
		4'd13: n_loc_oh_reg[85] = {2'd0, dist_reg[170], 13'd0};
		4'd14: n_loc_oh_reg[85] = {1'd0, dist_reg[170], 14'd0};
		4'd15: n_loc_oh_reg[85] = {dist_reg[170], 15'd0};
	endcase
	case(loc_reg[86])
		4'd0: n_loc_oh_reg[86] = {15'd0, dist_reg[169]};
		4'd1: n_loc_oh_reg[86] = {14'd0, dist_reg[169], 1'd0};
		4'd2: n_loc_oh_reg[86] = {13'd0, dist_reg[169], 2'd0};
		4'd3: n_loc_oh_reg[86] = {12'd0, dist_reg[169], 3'd0};
		4'd4: n_loc_oh_reg[86] = {11'd0, dist_reg[169], 4'd0};
		4'd5: n_loc_oh_reg[86] = {10'd0, dist_reg[169], 5'd0};
		4'd6: n_loc_oh_reg[86] = {9'd0, dist_reg[169], 6'd0};
		4'd7: n_loc_oh_reg[86] = {8'd0, dist_reg[169], 7'd0};
		4'd8: n_loc_oh_reg[86] = {7'd0, dist_reg[169], 8'd0};
		4'd9: n_loc_oh_reg[86] = {6'd0, dist_reg[169], 9'd0};
		4'd10: n_loc_oh_reg[86] = {5'd0, dist_reg[169], 10'd0};
		4'd11: n_loc_oh_reg[86] = {4'd0, dist_reg[169], 11'd0};
		4'd12: n_loc_oh_reg[86] = {3'd0, dist_reg[169], 12'd0};
		4'd13: n_loc_oh_reg[86] = {2'd0, dist_reg[169], 13'd0};
		4'd14: n_loc_oh_reg[86] = {1'd0, dist_reg[169], 14'd0};
		4'd15: n_loc_oh_reg[86] = {dist_reg[169], 15'd0};
	endcase
	case(loc_reg[87])
		4'd0: n_loc_oh_reg[87] = {15'd0, dist_reg[168]};
		4'd1: n_loc_oh_reg[87] = {14'd0, dist_reg[168], 1'd0};
		4'd2: n_loc_oh_reg[87] = {13'd0, dist_reg[168], 2'd0};
		4'd3: n_loc_oh_reg[87] = {12'd0, dist_reg[168], 3'd0};
		4'd4: n_loc_oh_reg[87] = {11'd0, dist_reg[168], 4'd0};
		4'd5: n_loc_oh_reg[87] = {10'd0, dist_reg[168], 5'd0};
		4'd6: n_loc_oh_reg[87] = {9'd0, dist_reg[168], 6'd0};
		4'd7: n_loc_oh_reg[87] = {8'd0, dist_reg[168], 7'd0};
		4'd8: n_loc_oh_reg[87] = {7'd0, dist_reg[168], 8'd0};
		4'd9: n_loc_oh_reg[87] = {6'd0, dist_reg[168], 9'd0};
		4'd10: n_loc_oh_reg[87] = {5'd0, dist_reg[168], 10'd0};
		4'd11: n_loc_oh_reg[87] = {4'd0, dist_reg[168], 11'd0};
		4'd12: n_loc_oh_reg[87] = {3'd0, dist_reg[168], 12'd0};
		4'd13: n_loc_oh_reg[87] = {2'd0, dist_reg[168], 13'd0};
		4'd14: n_loc_oh_reg[87] = {1'd0, dist_reg[168], 14'd0};
		4'd15: n_loc_oh_reg[87] = {dist_reg[168], 15'd0};
	endcase
	case(loc_reg[88])
		4'd0: n_loc_oh_reg[88] = {15'd0, dist_reg[167]};
		4'd1: n_loc_oh_reg[88] = {14'd0, dist_reg[167], 1'd0};
		4'd2: n_loc_oh_reg[88] = {13'd0, dist_reg[167], 2'd0};
		4'd3: n_loc_oh_reg[88] = {12'd0, dist_reg[167], 3'd0};
		4'd4: n_loc_oh_reg[88] = {11'd0, dist_reg[167], 4'd0};
		4'd5: n_loc_oh_reg[88] = {10'd0, dist_reg[167], 5'd0};
		4'd6: n_loc_oh_reg[88] = {9'd0, dist_reg[167], 6'd0};
		4'd7: n_loc_oh_reg[88] = {8'd0, dist_reg[167], 7'd0};
		4'd8: n_loc_oh_reg[88] = {7'd0, dist_reg[167], 8'd0};
		4'd9: n_loc_oh_reg[88] = {6'd0, dist_reg[167], 9'd0};
		4'd10: n_loc_oh_reg[88] = {5'd0, dist_reg[167], 10'd0};
		4'd11: n_loc_oh_reg[88] = {4'd0, dist_reg[167], 11'd0};
		4'd12: n_loc_oh_reg[88] = {3'd0, dist_reg[167], 12'd0};
		4'd13: n_loc_oh_reg[88] = {2'd0, dist_reg[167], 13'd0};
		4'd14: n_loc_oh_reg[88] = {1'd0, dist_reg[167], 14'd0};
		4'd15: n_loc_oh_reg[88] = {dist_reg[167], 15'd0};
	endcase
	case(loc_reg[89])
		4'd0: n_loc_oh_reg[89] = {15'd0, dist_reg[166]};
		4'd1: n_loc_oh_reg[89] = {14'd0, dist_reg[166], 1'd0};
		4'd2: n_loc_oh_reg[89] = {13'd0, dist_reg[166], 2'd0};
		4'd3: n_loc_oh_reg[89] = {12'd0, dist_reg[166], 3'd0};
		4'd4: n_loc_oh_reg[89] = {11'd0, dist_reg[166], 4'd0};
		4'd5: n_loc_oh_reg[89] = {10'd0, dist_reg[166], 5'd0};
		4'd6: n_loc_oh_reg[89] = {9'd0, dist_reg[166], 6'd0};
		4'd7: n_loc_oh_reg[89] = {8'd0, dist_reg[166], 7'd0};
		4'd8: n_loc_oh_reg[89] = {7'd0, dist_reg[166], 8'd0};
		4'd9: n_loc_oh_reg[89] = {6'd0, dist_reg[166], 9'd0};
		4'd10: n_loc_oh_reg[89] = {5'd0, dist_reg[166], 10'd0};
		4'd11: n_loc_oh_reg[89] = {4'd0, dist_reg[166], 11'd0};
		4'd12: n_loc_oh_reg[89] = {3'd0, dist_reg[166], 12'd0};
		4'd13: n_loc_oh_reg[89] = {2'd0, dist_reg[166], 13'd0};
		4'd14: n_loc_oh_reg[89] = {1'd0, dist_reg[166], 14'd0};
		4'd15: n_loc_oh_reg[89] = {dist_reg[166], 15'd0};
	endcase
	case(loc_reg[90])
		4'd0: n_loc_oh_reg[90] = {15'd0, dist_reg[165]};
		4'd1: n_loc_oh_reg[90] = {14'd0, dist_reg[165], 1'd0};
		4'd2: n_loc_oh_reg[90] = {13'd0, dist_reg[165], 2'd0};
		4'd3: n_loc_oh_reg[90] = {12'd0, dist_reg[165], 3'd0};
		4'd4: n_loc_oh_reg[90] = {11'd0, dist_reg[165], 4'd0};
		4'd5: n_loc_oh_reg[90] = {10'd0, dist_reg[165], 5'd0};
		4'd6: n_loc_oh_reg[90] = {9'd0, dist_reg[165], 6'd0};
		4'd7: n_loc_oh_reg[90] = {8'd0, dist_reg[165], 7'd0};
		4'd8: n_loc_oh_reg[90] = {7'd0, dist_reg[165], 8'd0};
		4'd9: n_loc_oh_reg[90] = {6'd0, dist_reg[165], 9'd0};
		4'd10: n_loc_oh_reg[90] = {5'd0, dist_reg[165], 10'd0};
		4'd11: n_loc_oh_reg[90] = {4'd0, dist_reg[165], 11'd0};
		4'd12: n_loc_oh_reg[90] = {3'd0, dist_reg[165], 12'd0};
		4'd13: n_loc_oh_reg[90] = {2'd0, dist_reg[165], 13'd0};
		4'd14: n_loc_oh_reg[90] = {1'd0, dist_reg[165], 14'd0};
		4'd15: n_loc_oh_reg[90] = {dist_reg[165], 15'd0};
	endcase
	case(loc_reg[91])
		4'd0: n_loc_oh_reg[91] = {15'd0, dist_reg[164]};
		4'd1: n_loc_oh_reg[91] = {14'd0, dist_reg[164], 1'd0};
		4'd2: n_loc_oh_reg[91] = {13'd0, dist_reg[164], 2'd0};
		4'd3: n_loc_oh_reg[91] = {12'd0, dist_reg[164], 3'd0};
		4'd4: n_loc_oh_reg[91] = {11'd0, dist_reg[164], 4'd0};
		4'd5: n_loc_oh_reg[91] = {10'd0, dist_reg[164], 5'd0};
		4'd6: n_loc_oh_reg[91] = {9'd0, dist_reg[164], 6'd0};
		4'd7: n_loc_oh_reg[91] = {8'd0, dist_reg[164], 7'd0};
		4'd8: n_loc_oh_reg[91] = {7'd0, dist_reg[164], 8'd0};
		4'd9: n_loc_oh_reg[91] = {6'd0, dist_reg[164], 9'd0};
		4'd10: n_loc_oh_reg[91] = {5'd0, dist_reg[164], 10'd0};
		4'd11: n_loc_oh_reg[91] = {4'd0, dist_reg[164], 11'd0};
		4'd12: n_loc_oh_reg[91] = {3'd0, dist_reg[164], 12'd0};
		4'd13: n_loc_oh_reg[91] = {2'd0, dist_reg[164], 13'd0};
		4'd14: n_loc_oh_reg[91] = {1'd0, dist_reg[164], 14'd0};
		4'd15: n_loc_oh_reg[91] = {dist_reg[164], 15'd0};
	endcase
	case(loc_reg[92])
		4'd0: n_loc_oh_reg[92] = {15'd0, dist_reg[163]};
		4'd1: n_loc_oh_reg[92] = {14'd0, dist_reg[163], 1'd0};
		4'd2: n_loc_oh_reg[92] = {13'd0, dist_reg[163], 2'd0};
		4'd3: n_loc_oh_reg[92] = {12'd0, dist_reg[163], 3'd0};
		4'd4: n_loc_oh_reg[92] = {11'd0, dist_reg[163], 4'd0};
		4'd5: n_loc_oh_reg[92] = {10'd0, dist_reg[163], 5'd0};
		4'd6: n_loc_oh_reg[92] = {9'd0, dist_reg[163], 6'd0};
		4'd7: n_loc_oh_reg[92] = {8'd0, dist_reg[163], 7'd0};
		4'd8: n_loc_oh_reg[92] = {7'd0, dist_reg[163], 8'd0};
		4'd9: n_loc_oh_reg[92] = {6'd0, dist_reg[163], 9'd0};
		4'd10: n_loc_oh_reg[92] = {5'd0, dist_reg[163], 10'd0};
		4'd11: n_loc_oh_reg[92] = {4'd0, dist_reg[163], 11'd0};
		4'd12: n_loc_oh_reg[92] = {3'd0, dist_reg[163], 12'd0};
		4'd13: n_loc_oh_reg[92] = {2'd0, dist_reg[163], 13'd0};
		4'd14: n_loc_oh_reg[92] = {1'd0, dist_reg[163], 14'd0};
		4'd15: n_loc_oh_reg[92] = {dist_reg[163], 15'd0};
	endcase
	case(loc_reg[93])
		4'd0: n_loc_oh_reg[93] = {15'd0, dist_reg[162]};
		4'd1: n_loc_oh_reg[93] = {14'd0, dist_reg[162], 1'd0};
		4'd2: n_loc_oh_reg[93] = {13'd0, dist_reg[162], 2'd0};
		4'd3: n_loc_oh_reg[93] = {12'd0, dist_reg[162], 3'd0};
		4'd4: n_loc_oh_reg[93] = {11'd0, dist_reg[162], 4'd0};
		4'd5: n_loc_oh_reg[93] = {10'd0, dist_reg[162], 5'd0};
		4'd6: n_loc_oh_reg[93] = {9'd0, dist_reg[162], 6'd0};
		4'd7: n_loc_oh_reg[93] = {8'd0, dist_reg[162], 7'd0};
		4'd8: n_loc_oh_reg[93] = {7'd0, dist_reg[162], 8'd0};
		4'd9: n_loc_oh_reg[93] = {6'd0, dist_reg[162], 9'd0};
		4'd10: n_loc_oh_reg[93] = {5'd0, dist_reg[162], 10'd0};
		4'd11: n_loc_oh_reg[93] = {4'd0, dist_reg[162], 11'd0};
		4'd12: n_loc_oh_reg[93] = {3'd0, dist_reg[162], 12'd0};
		4'd13: n_loc_oh_reg[93] = {2'd0, dist_reg[162], 13'd0};
		4'd14: n_loc_oh_reg[93] = {1'd0, dist_reg[162], 14'd0};
		4'd15: n_loc_oh_reg[93] = {dist_reg[162], 15'd0};
	endcase
	case(loc_reg[94])
		4'd0: n_loc_oh_reg[94] = {15'd0, dist_reg[161]};
		4'd1: n_loc_oh_reg[94] = {14'd0, dist_reg[161], 1'd0};
		4'd2: n_loc_oh_reg[94] = {13'd0, dist_reg[161], 2'd0};
		4'd3: n_loc_oh_reg[94] = {12'd0, dist_reg[161], 3'd0};
		4'd4: n_loc_oh_reg[94] = {11'd0, dist_reg[161], 4'd0};
		4'd5: n_loc_oh_reg[94] = {10'd0, dist_reg[161], 5'd0};
		4'd6: n_loc_oh_reg[94] = {9'd0, dist_reg[161], 6'd0};
		4'd7: n_loc_oh_reg[94] = {8'd0, dist_reg[161], 7'd0};
		4'd8: n_loc_oh_reg[94] = {7'd0, dist_reg[161], 8'd0};
		4'd9: n_loc_oh_reg[94] = {6'd0, dist_reg[161], 9'd0};
		4'd10: n_loc_oh_reg[94] = {5'd0, dist_reg[161], 10'd0};
		4'd11: n_loc_oh_reg[94] = {4'd0, dist_reg[161], 11'd0};
		4'd12: n_loc_oh_reg[94] = {3'd0, dist_reg[161], 12'd0};
		4'd13: n_loc_oh_reg[94] = {2'd0, dist_reg[161], 13'd0};
		4'd14: n_loc_oh_reg[94] = {1'd0, dist_reg[161], 14'd0};
		4'd15: n_loc_oh_reg[94] = {dist_reg[161], 15'd0};
	endcase
	case(loc_reg[95])
		4'd0: n_loc_oh_reg[95] = {15'd0, dist_reg[160]};
		4'd1: n_loc_oh_reg[95] = {14'd0, dist_reg[160], 1'd0};
		4'd2: n_loc_oh_reg[95] = {13'd0, dist_reg[160], 2'd0};
		4'd3: n_loc_oh_reg[95] = {12'd0, dist_reg[160], 3'd0};
		4'd4: n_loc_oh_reg[95] = {11'd0, dist_reg[160], 4'd0};
		4'd5: n_loc_oh_reg[95] = {10'd0, dist_reg[160], 5'd0};
		4'd6: n_loc_oh_reg[95] = {9'd0, dist_reg[160], 6'd0};
		4'd7: n_loc_oh_reg[95] = {8'd0, dist_reg[160], 7'd0};
		4'd8: n_loc_oh_reg[95] = {7'd0, dist_reg[160], 8'd0};
		4'd9: n_loc_oh_reg[95] = {6'd0, dist_reg[160], 9'd0};
		4'd10: n_loc_oh_reg[95] = {5'd0, dist_reg[160], 10'd0};
		4'd11: n_loc_oh_reg[95] = {4'd0, dist_reg[160], 11'd0};
		4'd12: n_loc_oh_reg[95] = {3'd0, dist_reg[160], 12'd0};
		4'd13: n_loc_oh_reg[95] = {2'd0, dist_reg[160], 13'd0};
		4'd14: n_loc_oh_reg[95] = {1'd0, dist_reg[160], 14'd0};
		4'd15: n_loc_oh_reg[95] = {dist_reg[160], 15'd0};
	endcase
	case(loc_reg[96])
		4'd0: n_loc_oh_reg[96] = {15'd0, dist_reg[159]};
		4'd1: n_loc_oh_reg[96] = {14'd0, dist_reg[159], 1'd0};
		4'd2: n_loc_oh_reg[96] = {13'd0, dist_reg[159], 2'd0};
		4'd3: n_loc_oh_reg[96] = {12'd0, dist_reg[159], 3'd0};
		4'd4: n_loc_oh_reg[96] = {11'd0, dist_reg[159], 4'd0};
		4'd5: n_loc_oh_reg[96] = {10'd0, dist_reg[159], 5'd0};
		4'd6: n_loc_oh_reg[96] = {9'd0, dist_reg[159], 6'd0};
		4'd7: n_loc_oh_reg[96] = {8'd0, dist_reg[159], 7'd0};
		4'd8: n_loc_oh_reg[96] = {7'd0, dist_reg[159], 8'd0};
		4'd9: n_loc_oh_reg[96] = {6'd0, dist_reg[159], 9'd0};
		4'd10: n_loc_oh_reg[96] = {5'd0, dist_reg[159], 10'd0};
		4'd11: n_loc_oh_reg[96] = {4'd0, dist_reg[159], 11'd0};
		4'd12: n_loc_oh_reg[96] = {3'd0, dist_reg[159], 12'd0};
		4'd13: n_loc_oh_reg[96] = {2'd0, dist_reg[159], 13'd0};
		4'd14: n_loc_oh_reg[96] = {1'd0, dist_reg[159], 14'd0};
		4'd15: n_loc_oh_reg[96] = {dist_reg[159], 15'd0};
	endcase
	case(loc_reg[97])
		4'd0: n_loc_oh_reg[97] = {15'd0, dist_reg[158]};
		4'd1: n_loc_oh_reg[97] = {14'd0, dist_reg[158], 1'd0};
		4'd2: n_loc_oh_reg[97] = {13'd0, dist_reg[158], 2'd0};
		4'd3: n_loc_oh_reg[97] = {12'd0, dist_reg[158], 3'd0};
		4'd4: n_loc_oh_reg[97] = {11'd0, dist_reg[158], 4'd0};
		4'd5: n_loc_oh_reg[97] = {10'd0, dist_reg[158], 5'd0};
		4'd6: n_loc_oh_reg[97] = {9'd0, dist_reg[158], 6'd0};
		4'd7: n_loc_oh_reg[97] = {8'd0, dist_reg[158], 7'd0};
		4'd8: n_loc_oh_reg[97] = {7'd0, dist_reg[158], 8'd0};
		4'd9: n_loc_oh_reg[97] = {6'd0, dist_reg[158], 9'd0};
		4'd10: n_loc_oh_reg[97] = {5'd0, dist_reg[158], 10'd0};
		4'd11: n_loc_oh_reg[97] = {4'd0, dist_reg[158], 11'd0};
		4'd12: n_loc_oh_reg[97] = {3'd0, dist_reg[158], 12'd0};
		4'd13: n_loc_oh_reg[97] = {2'd0, dist_reg[158], 13'd0};
		4'd14: n_loc_oh_reg[97] = {1'd0, dist_reg[158], 14'd0};
		4'd15: n_loc_oh_reg[97] = {dist_reg[158], 15'd0};
	endcase
	case(loc_reg[98])
		4'd0: n_loc_oh_reg[98] = {15'd0, dist_reg[157]};
		4'd1: n_loc_oh_reg[98] = {14'd0, dist_reg[157], 1'd0};
		4'd2: n_loc_oh_reg[98] = {13'd0, dist_reg[157], 2'd0};
		4'd3: n_loc_oh_reg[98] = {12'd0, dist_reg[157], 3'd0};
		4'd4: n_loc_oh_reg[98] = {11'd0, dist_reg[157], 4'd0};
		4'd5: n_loc_oh_reg[98] = {10'd0, dist_reg[157], 5'd0};
		4'd6: n_loc_oh_reg[98] = {9'd0, dist_reg[157], 6'd0};
		4'd7: n_loc_oh_reg[98] = {8'd0, dist_reg[157], 7'd0};
		4'd8: n_loc_oh_reg[98] = {7'd0, dist_reg[157], 8'd0};
		4'd9: n_loc_oh_reg[98] = {6'd0, dist_reg[157], 9'd0};
		4'd10: n_loc_oh_reg[98] = {5'd0, dist_reg[157], 10'd0};
		4'd11: n_loc_oh_reg[98] = {4'd0, dist_reg[157], 11'd0};
		4'd12: n_loc_oh_reg[98] = {3'd0, dist_reg[157], 12'd0};
		4'd13: n_loc_oh_reg[98] = {2'd0, dist_reg[157], 13'd0};
		4'd14: n_loc_oh_reg[98] = {1'd0, dist_reg[157], 14'd0};
		4'd15: n_loc_oh_reg[98] = {dist_reg[157], 15'd0};
	endcase
	case(loc_reg[99])
		4'd0: n_loc_oh_reg[99] = {15'd0, dist_reg[156]};
		4'd1: n_loc_oh_reg[99] = {14'd0, dist_reg[156], 1'd0};
		4'd2: n_loc_oh_reg[99] = {13'd0, dist_reg[156], 2'd0};
		4'd3: n_loc_oh_reg[99] = {12'd0, dist_reg[156], 3'd0};
		4'd4: n_loc_oh_reg[99] = {11'd0, dist_reg[156], 4'd0};
		4'd5: n_loc_oh_reg[99] = {10'd0, dist_reg[156], 5'd0};
		4'd6: n_loc_oh_reg[99] = {9'd0, dist_reg[156], 6'd0};
		4'd7: n_loc_oh_reg[99] = {8'd0, dist_reg[156], 7'd0};
		4'd8: n_loc_oh_reg[99] = {7'd0, dist_reg[156], 8'd0};
		4'd9: n_loc_oh_reg[99] = {6'd0, dist_reg[156], 9'd0};
		4'd10: n_loc_oh_reg[99] = {5'd0, dist_reg[156], 10'd0};
		4'd11: n_loc_oh_reg[99] = {4'd0, dist_reg[156], 11'd0};
		4'd12: n_loc_oh_reg[99] = {3'd0, dist_reg[156], 12'd0};
		4'd13: n_loc_oh_reg[99] = {2'd0, dist_reg[156], 13'd0};
		4'd14: n_loc_oh_reg[99] = {1'd0, dist_reg[156], 14'd0};
		4'd15: n_loc_oh_reg[99] = {dist_reg[156], 15'd0};
	endcase
	case(loc_reg[100])
		4'd0: n_loc_oh_reg[100] = {15'd0, dist_reg[155]};
		4'd1: n_loc_oh_reg[100] = {14'd0, dist_reg[155], 1'd0};
		4'd2: n_loc_oh_reg[100] = {13'd0, dist_reg[155], 2'd0};
		4'd3: n_loc_oh_reg[100] = {12'd0, dist_reg[155], 3'd0};
		4'd4: n_loc_oh_reg[100] = {11'd0, dist_reg[155], 4'd0};
		4'd5: n_loc_oh_reg[100] = {10'd0, dist_reg[155], 5'd0};
		4'd6: n_loc_oh_reg[100] = {9'd0, dist_reg[155], 6'd0};
		4'd7: n_loc_oh_reg[100] = {8'd0, dist_reg[155], 7'd0};
		4'd8: n_loc_oh_reg[100] = {7'd0, dist_reg[155], 8'd0};
		4'd9: n_loc_oh_reg[100] = {6'd0, dist_reg[155], 9'd0};
		4'd10: n_loc_oh_reg[100] = {5'd0, dist_reg[155], 10'd0};
		4'd11: n_loc_oh_reg[100] = {4'd0, dist_reg[155], 11'd0};
		4'd12: n_loc_oh_reg[100] = {3'd0, dist_reg[155], 12'd0};
		4'd13: n_loc_oh_reg[100] = {2'd0, dist_reg[155], 13'd0};
		4'd14: n_loc_oh_reg[100] = {1'd0, dist_reg[155], 14'd0};
		4'd15: n_loc_oh_reg[100] = {dist_reg[155], 15'd0};
	endcase
	case(loc_reg[101])
		4'd0: n_loc_oh_reg[101] = {15'd0, dist_reg[154]};
		4'd1: n_loc_oh_reg[101] = {14'd0, dist_reg[154], 1'd0};
		4'd2: n_loc_oh_reg[101] = {13'd0, dist_reg[154], 2'd0};
		4'd3: n_loc_oh_reg[101] = {12'd0, dist_reg[154], 3'd0};
		4'd4: n_loc_oh_reg[101] = {11'd0, dist_reg[154], 4'd0};
		4'd5: n_loc_oh_reg[101] = {10'd0, dist_reg[154], 5'd0};
		4'd6: n_loc_oh_reg[101] = {9'd0, dist_reg[154], 6'd0};
		4'd7: n_loc_oh_reg[101] = {8'd0, dist_reg[154], 7'd0};
		4'd8: n_loc_oh_reg[101] = {7'd0, dist_reg[154], 8'd0};
		4'd9: n_loc_oh_reg[101] = {6'd0, dist_reg[154], 9'd0};
		4'd10: n_loc_oh_reg[101] = {5'd0, dist_reg[154], 10'd0};
		4'd11: n_loc_oh_reg[101] = {4'd0, dist_reg[154], 11'd0};
		4'd12: n_loc_oh_reg[101] = {3'd0, dist_reg[154], 12'd0};
		4'd13: n_loc_oh_reg[101] = {2'd0, dist_reg[154], 13'd0};
		4'd14: n_loc_oh_reg[101] = {1'd0, dist_reg[154], 14'd0};
		4'd15: n_loc_oh_reg[101] = {dist_reg[154], 15'd0};
	endcase
	case(loc_reg[102])
		4'd0: n_loc_oh_reg[102] = {15'd0, dist_reg[153]};
		4'd1: n_loc_oh_reg[102] = {14'd0, dist_reg[153], 1'd0};
		4'd2: n_loc_oh_reg[102] = {13'd0, dist_reg[153], 2'd0};
		4'd3: n_loc_oh_reg[102] = {12'd0, dist_reg[153], 3'd0};
		4'd4: n_loc_oh_reg[102] = {11'd0, dist_reg[153], 4'd0};
		4'd5: n_loc_oh_reg[102] = {10'd0, dist_reg[153], 5'd0};
		4'd6: n_loc_oh_reg[102] = {9'd0, dist_reg[153], 6'd0};
		4'd7: n_loc_oh_reg[102] = {8'd0, dist_reg[153], 7'd0};
		4'd8: n_loc_oh_reg[102] = {7'd0, dist_reg[153], 8'd0};
		4'd9: n_loc_oh_reg[102] = {6'd0, dist_reg[153], 9'd0};
		4'd10: n_loc_oh_reg[102] = {5'd0, dist_reg[153], 10'd0};
		4'd11: n_loc_oh_reg[102] = {4'd0, dist_reg[153], 11'd0};
		4'd12: n_loc_oh_reg[102] = {3'd0, dist_reg[153], 12'd0};
		4'd13: n_loc_oh_reg[102] = {2'd0, dist_reg[153], 13'd0};
		4'd14: n_loc_oh_reg[102] = {1'd0, dist_reg[153], 14'd0};
		4'd15: n_loc_oh_reg[102] = {dist_reg[153], 15'd0};
	endcase
	case(loc_reg[103])
		4'd0: n_loc_oh_reg[103] = {15'd0, dist_reg[152]};
		4'd1: n_loc_oh_reg[103] = {14'd0, dist_reg[152], 1'd0};
		4'd2: n_loc_oh_reg[103] = {13'd0, dist_reg[152], 2'd0};
		4'd3: n_loc_oh_reg[103] = {12'd0, dist_reg[152], 3'd0};
		4'd4: n_loc_oh_reg[103] = {11'd0, dist_reg[152], 4'd0};
		4'd5: n_loc_oh_reg[103] = {10'd0, dist_reg[152], 5'd0};
		4'd6: n_loc_oh_reg[103] = {9'd0, dist_reg[152], 6'd0};
		4'd7: n_loc_oh_reg[103] = {8'd0, dist_reg[152], 7'd0};
		4'd8: n_loc_oh_reg[103] = {7'd0, dist_reg[152], 8'd0};
		4'd9: n_loc_oh_reg[103] = {6'd0, dist_reg[152], 9'd0};
		4'd10: n_loc_oh_reg[103] = {5'd0, dist_reg[152], 10'd0};
		4'd11: n_loc_oh_reg[103] = {4'd0, dist_reg[152], 11'd0};
		4'd12: n_loc_oh_reg[103] = {3'd0, dist_reg[152], 12'd0};
		4'd13: n_loc_oh_reg[103] = {2'd0, dist_reg[152], 13'd0};
		4'd14: n_loc_oh_reg[103] = {1'd0, dist_reg[152], 14'd0};
		4'd15: n_loc_oh_reg[103] = {dist_reg[152], 15'd0};
	endcase
	case(loc_reg[104])
		4'd0: n_loc_oh_reg[104] = {15'd0, dist_reg[151]};
		4'd1: n_loc_oh_reg[104] = {14'd0, dist_reg[151], 1'd0};
		4'd2: n_loc_oh_reg[104] = {13'd0, dist_reg[151], 2'd0};
		4'd3: n_loc_oh_reg[104] = {12'd0, dist_reg[151], 3'd0};
		4'd4: n_loc_oh_reg[104] = {11'd0, dist_reg[151], 4'd0};
		4'd5: n_loc_oh_reg[104] = {10'd0, dist_reg[151], 5'd0};
		4'd6: n_loc_oh_reg[104] = {9'd0, dist_reg[151], 6'd0};
		4'd7: n_loc_oh_reg[104] = {8'd0, dist_reg[151], 7'd0};
		4'd8: n_loc_oh_reg[104] = {7'd0, dist_reg[151], 8'd0};
		4'd9: n_loc_oh_reg[104] = {6'd0, dist_reg[151], 9'd0};
		4'd10: n_loc_oh_reg[104] = {5'd0, dist_reg[151], 10'd0};
		4'd11: n_loc_oh_reg[104] = {4'd0, dist_reg[151], 11'd0};
		4'd12: n_loc_oh_reg[104] = {3'd0, dist_reg[151], 12'd0};
		4'd13: n_loc_oh_reg[104] = {2'd0, dist_reg[151], 13'd0};
		4'd14: n_loc_oh_reg[104] = {1'd0, dist_reg[151], 14'd0};
		4'd15: n_loc_oh_reg[104] = {dist_reg[151], 15'd0};
	endcase
	case(loc_reg[105])
		4'd0: n_loc_oh_reg[105] = {15'd0, dist_reg[150]};
		4'd1: n_loc_oh_reg[105] = {14'd0, dist_reg[150], 1'd0};
		4'd2: n_loc_oh_reg[105] = {13'd0, dist_reg[150], 2'd0};
		4'd3: n_loc_oh_reg[105] = {12'd0, dist_reg[150], 3'd0};
		4'd4: n_loc_oh_reg[105] = {11'd0, dist_reg[150], 4'd0};
		4'd5: n_loc_oh_reg[105] = {10'd0, dist_reg[150], 5'd0};
		4'd6: n_loc_oh_reg[105] = {9'd0, dist_reg[150], 6'd0};
		4'd7: n_loc_oh_reg[105] = {8'd0, dist_reg[150], 7'd0};
		4'd8: n_loc_oh_reg[105] = {7'd0, dist_reg[150], 8'd0};
		4'd9: n_loc_oh_reg[105] = {6'd0, dist_reg[150], 9'd0};
		4'd10: n_loc_oh_reg[105] = {5'd0, dist_reg[150], 10'd0};
		4'd11: n_loc_oh_reg[105] = {4'd0, dist_reg[150], 11'd0};
		4'd12: n_loc_oh_reg[105] = {3'd0, dist_reg[150], 12'd0};
		4'd13: n_loc_oh_reg[105] = {2'd0, dist_reg[150], 13'd0};
		4'd14: n_loc_oh_reg[105] = {1'd0, dist_reg[150], 14'd0};
		4'd15: n_loc_oh_reg[105] = {dist_reg[150], 15'd0};
	endcase
	case(loc_reg[106])
		4'd0: n_loc_oh_reg[106] = {15'd0, dist_reg[149]};
		4'd1: n_loc_oh_reg[106] = {14'd0, dist_reg[149], 1'd0};
		4'd2: n_loc_oh_reg[106] = {13'd0, dist_reg[149], 2'd0};
		4'd3: n_loc_oh_reg[106] = {12'd0, dist_reg[149], 3'd0};
		4'd4: n_loc_oh_reg[106] = {11'd0, dist_reg[149], 4'd0};
		4'd5: n_loc_oh_reg[106] = {10'd0, dist_reg[149], 5'd0};
		4'd6: n_loc_oh_reg[106] = {9'd0, dist_reg[149], 6'd0};
		4'd7: n_loc_oh_reg[106] = {8'd0, dist_reg[149], 7'd0};
		4'd8: n_loc_oh_reg[106] = {7'd0, dist_reg[149], 8'd0};
		4'd9: n_loc_oh_reg[106] = {6'd0, dist_reg[149], 9'd0};
		4'd10: n_loc_oh_reg[106] = {5'd0, dist_reg[149], 10'd0};
		4'd11: n_loc_oh_reg[106] = {4'd0, dist_reg[149], 11'd0};
		4'd12: n_loc_oh_reg[106] = {3'd0, dist_reg[149], 12'd0};
		4'd13: n_loc_oh_reg[106] = {2'd0, dist_reg[149], 13'd0};
		4'd14: n_loc_oh_reg[106] = {1'd0, dist_reg[149], 14'd0};
		4'd15: n_loc_oh_reg[106] = {dist_reg[149], 15'd0};
	endcase
	case(loc_reg[107])
		4'd0: n_loc_oh_reg[107] = {15'd0, dist_reg[148]};
		4'd1: n_loc_oh_reg[107] = {14'd0, dist_reg[148], 1'd0};
		4'd2: n_loc_oh_reg[107] = {13'd0, dist_reg[148], 2'd0};
		4'd3: n_loc_oh_reg[107] = {12'd0, dist_reg[148], 3'd0};
		4'd4: n_loc_oh_reg[107] = {11'd0, dist_reg[148], 4'd0};
		4'd5: n_loc_oh_reg[107] = {10'd0, dist_reg[148], 5'd0};
		4'd6: n_loc_oh_reg[107] = {9'd0, dist_reg[148], 6'd0};
		4'd7: n_loc_oh_reg[107] = {8'd0, dist_reg[148], 7'd0};
		4'd8: n_loc_oh_reg[107] = {7'd0, dist_reg[148], 8'd0};
		4'd9: n_loc_oh_reg[107] = {6'd0, dist_reg[148], 9'd0};
		4'd10: n_loc_oh_reg[107] = {5'd0, dist_reg[148], 10'd0};
		4'd11: n_loc_oh_reg[107] = {4'd0, dist_reg[148], 11'd0};
		4'd12: n_loc_oh_reg[107] = {3'd0, dist_reg[148], 12'd0};
		4'd13: n_loc_oh_reg[107] = {2'd0, dist_reg[148], 13'd0};
		4'd14: n_loc_oh_reg[107] = {1'd0, dist_reg[148], 14'd0};
		4'd15: n_loc_oh_reg[107] = {dist_reg[148], 15'd0};
	endcase
	case(loc_reg[108])
		4'd0: n_loc_oh_reg[108] = {15'd0, dist_reg[147]};
		4'd1: n_loc_oh_reg[108] = {14'd0, dist_reg[147], 1'd0};
		4'd2: n_loc_oh_reg[108] = {13'd0, dist_reg[147], 2'd0};
		4'd3: n_loc_oh_reg[108] = {12'd0, dist_reg[147], 3'd0};
		4'd4: n_loc_oh_reg[108] = {11'd0, dist_reg[147], 4'd0};
		4'd5: n_loc_oh_reg[108] = {10'd0, dist_reg[147], 5'd0};
		4'd6: n_loc_oh_reg[108] = {9'd0, dist_reg[147], 6'd0};
		4'd7: n_loc_oh_reg[108] = {8'd0, dist_reg[147], 7'd0};
		4'd8: n_loc_oh_reg[108] = {7'd0, dist_reg[147], 8'd0};
		4'd9: n_loc_oh_reg[108] = {6'd0, dist_reg[147], 9'd0};
		4'd10: n_loc_oh_reg[108] = {5'd0, dist_reg[147], 10'd0};
		4'd11: n_loc_oh_reg[108] = {4'd0, dist_reg[147], 11'd0};
		4'd12: n_loc_oh_reg[108] = {3'd0, dist_reg[147], 12'd0};
		4'd13: n_loc_oh_reg[108] = {2'd0, dist_reg[147], 13'd0};
		4'd14: n_loc_oh_reg[108] = {1'd0, dist_reg[147], 14'd0};
		4'd15: n_loc_oh_reg[108] = {dist_reg[147], 15'd0};
	endcase
	case(loc_reg[109])
		4'd0: n_loc_oh_reg[109] = {15'd0, dist_reg[146]};
		4'd1: n_loc_oh_reg[109] = {14'd0, dist_reg[146], 1'd0};
		4'd2: n_loc_oh_reg[109] = {13'd0, dist_reg[146], 2'd0};
		4'd3: n_loc_oh_reg[109] = {12'd0, dist_reg[146], 3'd0};
		4'd4: n_loc_oh_reg[109] = {11'd0, dist_reg[146], 4'd0};
		4'd5: n_loc_oh_reg[109] = {10'd0, dist_reg[146], 5'd0};
		4'd6: n_loc_oh_reg[109] = {9'd0, dist_reg[146], 6'd0};
		4'd7: n_loc_oh_reg[109] = {8'd0, dist_reg[146], 7'd0};
		4'd8: n_loc_oh_reg[109] = {7'd0, dist_reg[146], 8'd0};
		4'd9: n_loc_oh_reg[109] = {6'd0, dist_reg[146], 9'd0};
		4'd10: n_loc_oh_reg[109] = {5'd0, dist_reg[146], 10'd0};
		4'd11: n_loc_oh_reg[109] = {4'd0, dist_reg[146], 11'd0};
		4'd12: n_loc_oh_reg[109] = {3'd0, dist_reg[146], 12'd0};
		4'd13: n_loc_oh_reg[109] = {2'd0, dist_reg[146], 13'd0};
		4'd14: n_loc_oh_reg[109] = {1'd0, dist_reg[146], 14'd0};
		4'd15: n_loc_oh_reg[109] = {dist_reg[146], 15'd0};
	endcase
	case(loc_reg[110])
		4'd0: n_loc_oh_reg[110] = {15'd0, dist_reg[145]};
		4'd1: n_loc_oh_reg[110] = {14'd0, dist_reg[145], 1'd0};
		4'd2: n_loc_oh_reg[110] = {13'd0, dist_reg[145], 2'd0};
		4'd3: n_loc_oh_reg[110] = {12'd0, dist_reg[145], 3'd0};
		4'd4: n_loc_oh_reg[110] = {11'd0, dist_reg[145], 4'd0};
		4'd5: n_loc_oh_reg[110] = {10'd0, dist_reg[145], 5'd0};
		4'd6: n_loc_oh_reg[110] = {9'd0, dist_reg[145], 6'd0};
		4'd7: n_loc_oh_reg[110] = {8'd0, dist_reg[145], 7'd0};
		4'd8: n_loc_oh_reg[110] = {7'd0, dist_reg[145], 8'd0};
		4'd9: n_loc_oh_reg[110] = {6'd0, dist_reg[145], 9'd0};
		4'd10: n_loc_oh_reg[110] = {5'd0, dist_reg[145], 10'd0};
		4'd11: n_loc_oh_reg[110] = {4'd0, dist_reg[145], 11'd0};
		4'd12: n_loc_oh_reg[110] = {3'd0, dist_reg[145], 12'd0};
		4'd13: n_loc_oh_reg[110] = {2'd0, dist_reg[145], 13'd0};
		4'd14: n_loc_oh_reg[110] = {1'd0, dist_reg[145], 14'd0};
		4'd15: n_loc_oh_reg[110] = {dist_reg[145], 15'd0};
	endcase
	case(loc_reg[111])
		4'd0: n_loc_oh_reg[111] = {15'd0, dist_reg[144]};
		4'd1: n_loc_oh_reg[111] = {14'd0, dist_reg[144], 1'd0};
		4'd2: n_loc_oh_reg[111] = {13'd0, dist_reg[144], 2'd0};
		4'd3: n_loc_oh_reg[111] = {12'd0, dist_reg[144], 3'd0};
		4'd4: n_loc_oh_reg[111] = {11'd0, dist_reg[144], 4'd0};
		4'd5: n_loc_oh_reg[111] = {10'd0, dist_reg[144], 5'd0};
		4'd6: n_loc_oh_reg[111] = {9'd0, dist_reg[144], 6'd0};
		4'd7: n_loc_oh_reg[111] = {8'd0, dist_reg[144], 7'd0};
		4'd8: n_loc_oh_reg[111] = {7'd0, dist_reg[144], 8'd0};
		4'd9: n_loc_oh_reg[111] = {6'd0, dist_reg[144], 9'd0};
		4'd10: n_loc_oh_reg[111] = {5'd0, dist_reg[144], 10'd0};
		4'd11: n_loc_oh_reg[111] = {4'd0, dist_reg[144], 11'd0};
		4'd12: n_loc_oh_reg[111] = {3'd0, dist_reg[144], 12'd0};
		4'd13: n_loc_oh_reg[111] = {2'd0, dist_reg[144], 13'd0};
		4'd14: n_loc_oh_reg[111] = {1'd0, dist_reg[144], 14'd0};
		4'd15: n_loc_oh_reg[111] = {dist_reg[144], 15'd0};
	endcase
	case(loc_reg[112])
		4'd0: n_loc_oh_reg[112] = {15'd0, dist_reg[143]};
		4'd1: n_loc_oh_reg[112] = {14'd0, dist_reg[143], 1'd0};
		4'd2: n_loc_oh_reg[112] = {13'd0, dist_reg[143], 2'd0};
		4'd3: n_loc_oh_reg[112] = {12'd0, dist_reg[143], 3'd0};
		4'd4: n_loc_oh_reg[112] = {11'd0, dist_reg[143], 4'd0};
		4'd5: n_loc_oh_reg[112] = {10'd0, dist_reg[143], 5'd0};
		4'd6: n_loc_oh_reg[112] = {9'd0, dist_reg[143], 6'd0};
		4'd7: n_loc_oh_reg[112] = {8'd0, dist_reg[143], 7'd0};
		4'd8: n_loc_oh_reg[112] = {7'd0, dist_reg[143], 8'd0};
		4'd9: n_loc_oh_reg[112] = {6'd0, dist_reg[143], 9'd0};
		4'd10: n_loc_oh_reg[112] = {5'd0, dist_reg[143], 10'd0};
		4'd11: n_loc_oh_reg[112] = {4'd0, dist_reg[143], 11'd0};
		4'd12: n_loc_oh_reg[112] = {3'd0, dist_reg[143], 12'd0};
		4'd13: n_loc_oh_reg[112] = {2'd0, dist_reg[143], 13'd0};
		4'd14: n_loc_oh_reg[112] = {1'd0, dist_reg[143], 14'd0};
		4'd15: n_loc_oh_reg[112] = {dist_reg[143], 15'd0};
	endcase
	case(loc_reg[113])
		4'd0: n_loc_oh_reg[113] = {15'd0, dist_reg[142]};
		4'd1: n_loc_oh_reg[113] = {14'd0, dist_reg[142], 1'd0};
		4'd2: n_loc_oh_reg[113] = {13'd0, dist_reg[142], 2'd0};
		4'd3: n_loc_oh_reg[113] = {12'd0, dist_reg[142], 3'd0};
		4'd4: n_loc_oh_reg[113] = {11'd0, dist_reg[142], 4'd0};
		4'd5: n_loc_oh_reg[113] = {10'd0, dist_reg[142], 5'd0};
		4'd6: n_loc_oh_reg[113] = {9'd0, dist_reg[142], 6'd0};
		4'd7: n_loc_oh_reg[113] = {8'd0, dist_reg[142], 7'd0};
		4'd8: n_loc_oh_reg[113] = {7'd0, dist_reg[142], 8'd0};
		4'd9: n_loc_oh_reg[113] = {6'd0, dist_reg[142], 9'd0};
		4'd10: n_loc_oh_reg[113] = {5'd0, dist_reg[142], 10'd0};
		4'd11: n_loc_oh_reg[113] = {4'd0, dist_reg[142], 11'd0};
		4'd12: n_loc_oh_reg[113] = {3'd0, dist_reg[142], 12'd0};
		4'd13: n_loc_oh_reg[113] = {2'd0, dist_reg[142], 13'd0};
		4'd14: n_loc_oh_reg[113] = {1'd0, dist_reg[142], 14'd0};
		4'd15: n_loc_oh_reg[113] = {dist_reg[142], 15'd0};
	endcase
	case(loc_reg[114])
		4'd0: n_loc_oh_reg[114] = {15'd0, dist_reg[141]};
		4'd1: n_loc_oh_reg[114] = {14'd0, dist_reg[141], 1'd0};
		4'd2: n_loc_oh_reg[114] = {13'd0, dist_reg[141], 2'd0};
		4'd3: n_loc_oh_reg[114] = {12'd0, dist_reg[141], 3'd0};
		4'd4: n_loc_oh_reg[114] = {11'd0, dist_reg[141], 4'd0};
		4'd5: n_loc_oh_reg[114] = {10'd0, dist_reg[141], 5'd0};
		4'd6: n_loc_oh_reg[114] = {9'd0, dist_reg[141], 6'd0};
		4'd7: n_loc_oh_reg[114] = {8'd0, dist_reg[141], 7'd0};
		4'd8: n_loc_oh_reg[114] = {7'd0, dist_reg[141], 8'd0};
		4'd9: n_loc_oh_reg[114] = {6'd0, dist_reg[141], 9'd0};
		4'd10: n_loc_oh_reg[114] = {5'd0, dist_reg[141], 10'd0};
		4'd11: n_loc_oh_reg[114] = {4'd0, dist_reg[141], 11'd0};
		4'd12: n_loc_oh_reg[114] = {3'd0, dist_reg[141], 12'd0};
		4'd13: n_loc_oh_reg[114] = {2'd0, dist_reg[141], 13'd0};
		4'd14: n_loc_oh_reg[114] = {1'd0, dist_reg[141], 14'd0};
		4'd15: n_loc_oh_reg[114] = {dist_reg[141], 15'd0};
	endcase
	case(loc_reg[115])
		4'd0: n_loc_oh_reg[115] = {15'd0, dist_reg[140]};
		4'd1: n_loc_oh_reg[115] = {14'd0, dist_reg[140], 1'd0};
		4'd2: n_loc_oh_reg[115] = {13'd0, dist_reg[140], 2'd0};
		4'd3: n_loc_oh_reg[115] = {12'd0, dist_reg[140], 3'd0};
		4'd4: n_loc_oh_reg[115] = {11'd0, dist_reg[140], 4'd0};
		4'd5: n_loc_oh_reg[115] = {10'd0, dist_reg[140], 5'd0};
		4'd6: n_loc_oh_reg[115] = {9'd0, dist_reg[140], 6'd0};
		4'd7: n_loc_oh_reg[115] = {8'd0, dist_reg[140], 7'd0};
		4'd8: n_loc_oh_reg[115] = {7'd0, dist_reg[140], 8'd0};
		4'd9: n_loc_oh_reg[115] = {6'd0, dist_reg[140], 9'd0};
		4'd10: n_loc_oh_reg[115] = {5'd0, dist_reg[140], 10'd0};
		4'd11: n_loc_oh_reg[115] = {4'd0, dist_reg[140], 11'd0};
		4'd12: n_loc_oh_reg[115] = {3'd0, dist_reg[140], 12'd0};
		4'd13: n_loc_oh_reg[115] = {2'd0, dist_reg[140], 13'd0};
		4'd14: n_loc_oh_reg[115] = {1'd0, dist_reg[140], 14'd0};
		4'd15: n_loc_oh_reg[115] = {dist_reg[140], 15'd0};
	endcase
	case(loc_reg[116])
		4'd0: n_loc_oh_reg[116] = {15'd0, dist_reg[139]};
		4'd1: n_loc_oh_reg[116] = {14'd0, dist_reg[139], 1'd0};
		4'd2: n_loc_oh_reg[116] = {13'd0, dist_reg[139], 2'd0};
		4'd3: n_loc_oh_reg[116] = {12'd0, dist_reg[139], 3'd0};
		4'd4: n_loc_oh_reg[116] = {11'd0, dist_reg[139], 4'd0};
		4'd5: n_loc_oh_reg[116] = {10'd0, dist_reg[139], 5'd0};
		4'd6: n_loc_oh_reg[116] = {9'd0, dist_reg[139], 6'd0};
		4'd7: n_loc_oh_reg[116] = {8'd0, dist_reg[139], 7'd0};
		4'd8: n_loc_oh_reg[116] = {7'd0, dist_reg[139], 8'd0};
		4'd9: n_loc_oh_reg[116] = {6'd0, dist_reg[139], 9'd0};
		4'd10: n_loc_oh_reg[116] = {5'd0, dist_reg[139], 10'd0};
		4'd11: n_loc_oh_reg[116] = {4'd0, dist_reg[139], 11'd0};
		4'd12: n_loc_oh_reg[116] = {3'd0, dist_reg[139], 12'd0};
		4'd13: n_loc_oh_reg[116] = {2'd0, dist_reg[139], 13'd0};
		4'd14: n_loc_oh_reg[116] = {1'd0, dist_reg[139], 14'd0};
		4'd15: n_loc_oh_reg[116] = {dist_reg[139], 15'd0};
	endcase
	case(loc_reg[117])
		4'd0: n_loc_oh_reg[117] = {15'd0, dist_reg[138]};
		4'd1: n_loc_oh_reg[117] = {14'd0, dist_reg[138], 1'd0};
		4'd2: n_loc_oh_reg[117] = {13'd0, dist_reg[138], 2'd0};
		4'd3: n_loc_oh_reg[117] = {12'd0, dist_reg[138], 3'd0};
		4'd4: n_loc_oh_reg[117] = {11'd0, dist_reg[138], 4'd0};
		4'd5: n_loc_oh_reg[117] = {10'd0, dist_reg[138], 5'd0};
		4'd6: n_loc_oh_reg[117] = {9'd0, dist_reg[138], 6'd0};
		4'd7: n_loc_oh_reg[117] = {8'd0, dist_reg[138], 7'd0};
		4'd8: n_loc_oh_reg[117] = {7'd0, dist_reg[138], 8'd0};
		4'd9: n_loc_oh_reg[117] = {6'd0, dist_reg[138], 9'd0};
		4'd10: n_loc_oh_reg[117] = {5'd0, dist_reg[138], 10'd0};
		4'd11: n_loc_oh_reg[117] = {4'd0, dist_reg[138], 11'd0};
		4'd12: n_loc_oh_reg[117] = {3'd0, dist_reg[138], 12'd0};
		4'd13: n_loc_oh_reg[117] = {2'd0, dist_reg[138], 13'd0};
		4'd14: n_loc_oh_reg[117] = {1'd0, dist_reg[138], 14'd0};
		4'd15: n_loc_oh_reg[117] = {dist_reg[138], 15'd0};
	endcase
	case(loc_reg[118])
		4'd0: n_loc_oh_reg[118] = {15'd0, dist_reg[137]};
		4'd1: n_loc_oh_reg[118] = {14'd0, dist_reg[137], 1'd0};
		4'd2: n_loc_oh_reg[118] = {13'd0, dist_reg[137], 2'd0};
		4'd3: n_loc_oh_reg[118] = {12'd0, dist_reg[137], 3'd0};
		4'd4: n_loc_oh_reg[118] = {11'd0, dist_reg[137], 4'd0};
		4'd5: n_loc_oh_reg[118] = {10'd0, dist_reg[137], 5'd0};
		4'd6: n_loc_oh_reg[118] = {9'd0, dist_reg[137], 6'd0};
		4'd7: n_loc_oh_reg[118] = {8'd0, dist_reg[137], 7'd0};
		4'd8: n_loc_oh_reg[118] = {7'd0, dist_reg[137], 8'd0};
		4'd9: n_loc_oh_reg[118] = {6'd0, dist_reg[137], 9'd0};
		4'd10: n_loc_oh_reg[118] = {5'd0, dist_reg[137], 10'd0};
		4'd11: n_loc_oh_reg[118] = {4'd0, dist_reg[137], 11'd0};
		4'd12: n_loc_oh_reg[118] = {3'd0, dist_reg[137], 12'd0};
		4'd13: n_loc_oh_reg[118] = {2'd0, dist_reg[137], 13'd0};
		4'd14: n_loc_oh_reg[118] = {1'd0, dist_reg[137], 14'd0};
		4'd15: n_loc_oh_reg[118] = {dist_reg[137], 15'd0};
	endcase
	case(loc_reg[119])
		4'd0: n_loc_oh_reg[119] = {15'd0, dist_reg[136]};
		4'd1: n_loc_oh_reg[119] = {14'd0, dist_reg[136], 1'd0};
		4'd2: n_loc_oh_reg[119] = {13'd0, dist_reg[136], 2'd0};
		4'd3: n_loc_oh_reg[119] = {12'd0, dist_reg[136], 3'd0};
		4'd4: n_loc_oh_reg[119] = {11'd0, dist_reg[136], 4'd0};
		4'd5: n_loc_oh_reg[119] = {10'd0, dist_reg[136], 5'd0};
		4'd6: n_loc_oh_reg[119] = {9'd0, dist_reg[136], 6'd0};
		4'd7: n_loc_oh_reg[119] = {8'd0, dist_reg[136], 7'd0};
		4'd8: n_loc_oh_reg[119] = {7'd0, dist_reg[136], 8'd0};
		4'd9: n_loc_oh_reg[119] = {6'd0, dist_reg[136], 9'd0};
		4'd10: n_loc_oh_reg[119] = {5'd0, dist_reg[136], 10'd0};
		4'd11: n_loc_oh_reg[119] = {4'd0, dist_reg[136], 11'd0};
		4'd12: n_loc_oh_reg[119] = {3'd0, dist_reg[136], 12'd0};
		4'd13: n_loc_oh_reg[119] = {2'd0, dist_reg[136], 13'd0};
		4'd14: n_loc_oh_reg[119] = {1'd0, dist_reg[136], 14'd0};
		4'd15: n_loc_oh_reg[119] = {dist_reg[136], 15'd0};
	endcase
	case(loc_reg[120])
		4'd0: n_loc_oh_reg[120] = {15'd0, dist_reg[135]};
		4'd1: n_loc_oh_reg[120] = {14'd0, dist_reg[135], 1'd0};
		4'd2: n_loc_oh_reg[120] = {13'd0, dist_reg[135], 2'd0};
		4'd3: n_loc_oh_reg[120] = {12'd0, dist_reg[135], 3'd0};
		4'd4: n_loc_oh_reg[120] = {11'd0, dist_reg[135], 4'd0};
		4'd5: n_loc_oh_reg[120] = {10'd0, dist_reg[135], 5'd0};
		4'd6: n_loc_oh_reg[120] = {9'd0, dist_reg[135], 6'd0};
		4'd7: n_loc_oh_reg[120] = {8'd0, dist_reg[135], 7'd0};
		4'd8: n_loc_oh_reg[120] = {7'd0, dist_reg[135], 8'd0};
		4'd9: n_loc_oh_reg[120] = {6'd0, dist_reg[135], 9'd0};
		4'd10: n_loc_oh_reg[120] = {5'd0, dist_reg[135], 10'd0};
		4'd11: n_loc_oh_reg[120] = {4'd0, dist_reg[135], 11'd0};
		4'd12: n_loc_oh_reg[120] = {3'd0, dist_reg[135], 12'd0};
		4'd13: n_loc_oh_reg[120] = {2'd0, dist_reg[135], 13'd0};
		4'd14: n_loc_oh_reg[120] = {1'd0, dist_reg[135], 14'd0};
		4'd15: n_loc_oh_reg[120] = {dist_reg[135], 15'd0};
	endcase
	case(loc_reg[121])
		4'd0: n_loc_oh_reg[121] = {15'd0, dist_reg[134]};
		4'd1: n_loc_oh_reg[121] = {14'd0, dist_reg[134], 1'd0};
		4'd2: n_loc_oh_reg[121] = {13'd0, dist_reg[134], 2'd0};
		4'd3: n_loc_oh_reg[121] = {12'd0, dist_reg[134], 3'd0};
		4'd4: n_loc_oh_reg[121] = {11'd0, dist_reg[134], 4'd0};
		4'd5: n_loc_oh_reg[121] = {10'd0, dist_reg[134], 5'd0};
		4'd6: n_loc_oh_reg[121] = {9'd0, dist_reg[134], 6'd0};
		4'd7: n_loc_oh_reg[121] = {8'd0, dist_reg[134], 7'd0};
		4'd8: n_loc_oh_reg[121] = {7'd0, dist_reg[134], 8'd0};
		4'd9: n_loc_oh_reg[121] = {6'd0, dist_reg[134], 9'd0};
		4'd10: n_loc_oh_reg[121] = {5'd0, dist_reg[134], 10'd0};
		4'd11: n_loc_oh_reg[121] = {4'd0, dist_reg[134], 11'd0};
		4'd12: n_loc_oh_reg[121] = {3'd0, dist_reg[134], 12'd0};
		4'd13: n_loc_oh_reg[121] = {2'd0, dist_reg[134], 13'd0};
		4'd14: n_loc_oh_reg[121] = {1'd0, dist_reg[134], 14'd0};
		4'd15: n_loc_oh_reg[121] = {dist_reg[134], 15'd0};
	endcase
	case(loc_reg[122])
		4'd0: n_loc_oh_reg[122] = {15'd0, dist_reg[133]};
		4'd1: n_loc_oh_reg[122] = {14'd0, dist_reg[133], 1'd0};
		4'd2: n_loc_oh_reg[122] = {13'd0, dist_reg[133], 2'd0};
		4'd3: n_loc_oh_reg[122] = {12'd0, dist_reg[133], 3'd0};
		4'd4: n_loc_oh_reg[122] = {11'd0, dist_reg[133], 4'd0};
		4'd5: n_loc_oh_reg[122] = {10'd0, dist_reg[133], 5'd0};
		4'd6: n_loc_oh_reg[122] = {9'd0, dist_reg[133], 6'd0};
		4'd7: n_loc_oh_reg[122] = {8'd0, dist_reg[133], 7'd0};
		4'd8: n_loc_oh_reg[122] = {7'd0, dist_reg[133], 8'd0};
		4'd9: n_loc_oh_reg[122] = {6'd0, dist_reg[133], 9'd0};
		4'd10: n_loc_oh_reg[122] = {5'd0, dist_reg[133], 10'd0};
		4'd11: n_loc_oh_reg[122] = {4'd0, dist_reg[133], 11'd0};
		4'd12: n_loc_oh_reg[122] = {3'd0, dist_reg[133], 12'd0};
		4'd13: n_loc_oh_reg[122] = {2'd0, dist_reg[133], 13'd0};
		4'd14: n_loc_oh_reg[122] = {1'd0, dist_reg[133], 14'd0};
		4'd15: n_loc_oh_reg[122] = {dist_reg[133], 15'd0};
	endcase
	case(loc_reg[123])
		4'd0: n_loc_oh_reg[123] = {15'd0, dist_reg[132]};
		4'd1: n_loc_oh_reg[123] = {14'd0, dist_reg[132], 1'd0};
		4'd2: n_loc_oh_reg[123] = {13'd0, dist_reg[132], 2'd0};
		4'd3: n_loc_oh_reg[123] = {12'd0, dist_reg[132], 3'd0};
		4'd4: n_loc_oh_reg[123] = {11'd0, dist_reg[132], 4'd0};
		4'd5: n_loc_oh_reg[123] = {10'd0, dist_reg[132], 5'd0};
		4'd6: n_loc_oh_reg[123] = {9'd0, dist_reg[132], 6'd0};
		4'd7: n_loc_oh_reg[123] = {8'd0, dist_reg[132], 7'd0};
		4'd8: n_loc_oh_reg[123] = {7'd0, dist_reg[132], 8'd0};
		4'd9: n_loc_oh_reg[123] = {6'd0, dist_reg[132], 9'd0};
		4'd10: n_loc_oh_reg[123] = {5'd0, dist_reg[132], 10'd0};
		4'd11: n_loc_oh_reg[123] = {4'd0, dist_reg[132], 11'd0};
		4'd12: n_loc_oh_reg[123] = {3'd0, dist_reg[132], 12'd0};
		4'd13: n_loc_oh_reg[123] = {2'd0, dist_reg[132], 13'd0};
		4'd14: n_loc_oh_reg[123] = {1'd0, dist_reg[132], 14'd0};
		4'd15: n_loc_oh_reg[123] = {dist_reg[132], 15'd0};
	endcase
	case(loc_reg[124])
		4'd0: n_loc_oh_reg[124] = {15'd0, dist_reg[131]};
		4'd1: n_loc_oh_reg[124] = {14'd0, dist_reg[131], 1'd0};
		4'd2: n_loc_oh_reg[124] = {13'd0, dist_reg[131], 2'd0};
		4'd3: n_loc_oh_reg[124] = {12'd0, dist_reg[131], 3'd0};
		4'd4: n_loc_oh_reg[124] = {11'd0, dist_reg[131], 4'd0};
		4'd5: n_loc_oh_reg[124] = {10'd0, dist_reg[131], 5'd0};
		4'd6: n_loc_oh_reg[124] = {9'd0, dist_reg[131], 6'd0};
		4'd7: n_loc_oh_reg[124] = {8'd0, dist_reg[131], 7'd0};
		4'd8: n_loc_oh_reg[124] = {7'd0, dist_reg[131], 8'd0};
		4'd9: n_loc_oh_reg[124] = {6'd0, dist_reg[131], 9'd0};
		4'd10: n_loc_oh_reg[124] = {5'd0, dist_reg[131], 10'd0};
		4'd11: n_loc_oh_reg[124] = {4'd0, dist_reg[131], 11'd0};
		4'd12: n_loc_oh_reg[124] = {3'd0, dist_reg[131], 12'd0};
		4'd13: n_loc_oh_reg[124] = {2'd0, dist_reg[131], 13'd0};
		4'd14: n_loc_oh_reg[124] = {1'd0, dist_reg[131], 14'd0};
		4'd15: n_loc_oh_reg[124] = {dist_reg[131], 15'd0};
	endcase
	case(loc_reg[125])
		4'd0: n_loc_oh_reg[125] = {15'd0, dist_reg[130]};
		4'd1: n_loc_oh_reg[125] = {14'd0, dist_reg[130], 1'd0};
		4'd2: n_loc_oh_reg[125] = {13'd0, dist_reg[130], 2'd0};
		4'd3: n_loc_oh_reg[125] = {12'd0, dist_reg[130], 3'd0};
		4'd4: n_loc_oh_reg[125] = {11'd0, dist_reg[130], 4'd0};
		4'd5: n_loc_oh_reg[125] = {10'd0, dist_reg[130], 5'd0};
		4'd6: n_loc_oh_reg[125] = {9'd0, dist_reg[130], 6'd0};
		4'd7: n_loc_oh_reg[125] = {8'd0, dist_reg[130], 7'd0};
		4'd8: n_loc_oh_reg[125] = {7'd0, dist_reg[130], 8'd0};
		4'd9: n_loc_oh_reg[125] = {6'd0, dist_reg[130], 9'd0};
		4'd10: n_loc_oh_reg[125] = {5'd0, dist_reg[130], 10'd0};
		4'd11: n_loc_oh_reg[125] = {4'd0, dist_reg[130], 11'd0};
		4'd12: n_loc_oh_reg[125] = {3'd0, dist_reg[130], 12'd0};
		4'd13: n_loc_oh_reg[125] = {2'd0, dist_reg[130], 13'd0};
		4'd14: n_loc_oh_reg[125] = {1'd0, dist_reg[130], 14'd0};
		4'd15: n_loc_oh_reg[125] = {dist_reg[130], 15'd0};
	endcase
	case(loc_reg[126])
		4'd0: n_loc_oh_reg[126] = {15'd0, dist_reg[129]};
		4'd1: n_loc_oh_reg[126] = {14'd0, dist_reg[129], 1'd0};
		4'd2: n_loc_oh_reg[126] = {13'd0, dist_reg[129], 2'd0};
		4'd3: n_loc_oh_reg[126] = {12'd0, dist_reg[129], 3'd0};
		4'd4: n_loc_oh_reg[126] = {11'd0, dist_reg[129], 4'd0};
		4'd5: n_loc_oh_reg[126] = {10'd0, dist_reg[129], 5'd0};
		4'd6: n_loc_oh_reg[126] = {9'd0, dist_reg[129], 6'd0};
		4'd7: n_loc_oh_reg[126] = {8'd0, dist_reg[129], 7'd0};
		4'd8: n_loc_oh_reg[126] = {7'd0, dist_reg[129], 8'd0};
		4'd9: n_loc_oh_reg[126] = {6'd0, dist_reg[129], 9'd0};
		4'd10: n_loc_oh_reg[126] = {5'd0, dist_reg[129], 10'd0};
		4'd11: n_loc_oh_reg[126] = {4'd0, dist_reg[129], 11'd0};
		4'd12: n_loc_oh_reg[126] = {3'd0, dist_reg[129], 12'd0};
		4'd13: n_loc_oh_reg[126] = {2'd0, dist_reg[129], 13'd0};
		4'd14: n_loc_oh_reg[126] = {1'd0, dist_reg[129], 14'd0};
		4'd15: n_loc_oh_reg[126] = {dist_reg[129], 15'd0};
	endcase
	case(loc_reg[127])
		4'd0: n_loc_oh_reg[127] = {15'd0, dist_reg[128]};
		4'd1: n_loc_oh_reg[127] = {14'd0, dist_reg[128], 1'd0};
		4'd2: n_loc_oh_reg[127] = {13'd0, dist_reg[128], 2'd0};
		4'd3: n_loc_oh_reg[127] = {12'd0, dist_reg[128], 3'd0};
		4'd4: n_loc_oh_reg[127] = {11'd0, dist_reg[128], 4'd0};
		4'd5: n_loc_oh_reg[127] = {10'd0, dist_reg[128], 5'd0};
		4'd6: n_loc_oh_reg[127] = {9'd0, dist_reg[128], 6'd0};
		4'd7: n_loc_oh_reg[127] = {8'd0, dist_reg[128], 7'd0};
		4'd8: n_loc_oh_reg[127] = {7'd0, dist_reg[128], 8'd0};
		4'd9: n_loc_oh_reg[127] = {6'd0, dist_reg[128], 9'd0};
		4'd10: n_loc_oh_reg[127] = {5'd0, dist_reg[128], 10'd0};
		4'd11: n_loc_oh_reg[127] = {4'd0, dist_reg[128], 11'd0};
		4'd12: n_loc_oh_reg[127] = {3'd0, dist_reg[128], 12'd0};
		4'd13: n_loc_oh_reg[127] = {2'd0, dist_reg[128], 13'd0};
		4'd14: n_loc_oh_reg[127] = {1'd0, dist_reg[128], 14'd0};
		4'd15: n_loc_oh_reg[127] = {dist_reg[128], 15'd0};
	endcase
	case(loc_reg[128])
		4'd0: n_loc_oh_reg[128] = {15'd0, dist_reg[127]};
		4'd1: n_loc_oh_reg[128] = {14'd0, dist_reg[127], 1'd0};
		4'd2: n_loc_oh_reg[128] = {13'd0, dist_reg[127], 2'd0};
		4'd3: n_loc_oh_reg[128] = {12'd0, dist_reg[127], 3'd0};
		4'd4: n_loc_oh_reg[128] = {11'd0, dist_reg[127], 4'd0};
		4'd5: n_loc_oh_reg[128] = {10'd0, dist_reg[127], 5'd0};
		4'd6: n_loc_oh_reg[128] = {9'd0, dist_reg[127], 6'd0};
		4'd7: n_loc_oh_reg[128] = {8'd0, dist_reg[127], 7'd0};
		4'd8: n_loc_oh_reg[128] = {7'd0, dist_reg[127], 8'd0};
		4'd9: n_loc_oh_reg[128] = {6'd0, dist_reg[127], 9'd0};
		4'd10: n_loc_oh_reg[128] = {5'd0, dist_reg[127], 10'd0};
		4'd11: n_loc_oh_reg[128] = {4'd0, dist_reg[127], 11'd0};
		4'd12: n_loc_oh_reg[128] = {3'd0, dist_reg[127], 12'd0};
		4'd13: n_loc_oh_reg[128] = {2'd0, dist_reg[127], 13'd0};
		4'd14: n_loc_oh_reg[128] = {1'd0, dist_reg[127], 14'd0};
		4'd15: n_loc_oh_reg[128] = {dist_reg[127], 15'd0};
	endcase
	case(loc_reg[129])
		4'd0: n_loc_oh_reg[129] = {15'd0, dist_reg[126]};
		4'd1: n_loc_oh_reg[129] = {14'd0, dist_reg[126], 1'd0};
		4'd2: n_loc_oh_reg[129] = {13'd0, dist_reg[126], 2'd0};
		4'd3: n_loc_oh_reg[129] = {12'd0, dist_reg[126], 3'd0};
		4'd4: n_loc_oh_reg[129] = {11'd0, dist_reg[126], 4'd0};
		4'd5: n_loc_oh_reg[129] = {10'd0, dist_reg[126], 5'd0};
		4'd6: n_loc_oh_reg[129] = {9'd0, dist_reg[126], 6'd0};
		4'd7: n_loc_oh_reg[129] = {8'd0, dist_reg[126], 7'd0};
		4'd8: n_loc_oh_reg[129] = {7'd0, dist_reg[126], 8'd0};
		4'd9: n_loc_oh_reg[129] = {6'd0, dist_reg[126], 9'd0};
		4'd10: n_loc_oh_reg[129] = {5'd0, dist_reg[126], 10'd0};
		4'd11: n_loc_oh_reg[129] = {4'd0, dist_reg[126], 11'd0};
		4'd12: n_loc_oh_reg[129] = {3'd0, dist_reg[126], 12'd0};
		4'd13: n_loc_oh_reg[129] = {2'd0, dist_reg[126], 13'd0};
		4'd14: n_loc_oh_reg[129] = {1'd0, dist_reg[126], 14'd0};
		4'd15: n_loc_oh_reg[129] = {dist_reg[126], 15'd0};
	endcase
	case(loc_reg[130])
		4'd0: n_loc_oh_reg[130] = {15'd0, dist_reg[125]};
		4'd1: n_loc_oh_reg[130] = {14'd0, dist_reg[125], 1'd0};
		4'd2: n_loc_oh_reg[130] = {13'd0, dist_reg[125], 2'd0};
		4'd3: n_loc_oh_reg[130] = {12'd0, dist_reg[125], 3'd0};
		4'd4: n_loc_oh_reg[130] = {11'd0, dist_reg[125], 4'd0};
		4'd5: n_loc_oh_reg[130] = {10'd0, dist_reg[125], 5'd0};
		4'd6: n_loc_oh_reg[130] = {9'd0, dist_reg[125], 6'd0};
		4'd7: n_loc_oh_reg[130] = {8'd0, dist_reg[125], 7'd0};
		4'd8: n_loc_oh_reg[130] = {7'd0, dist_reg[125], 8'd0};
		4'd9: n_loc_oh_reg[130] = {6'd0, dist_reg[125], 9'd0};
		4'd10: n_loc_oh_reg[130] = {5'd0, dist_reg[125], 10'd0};
		4'd11: n_loc_oh_reg[130] = {4'd0, dist_reg[125], 11'd0};
		4'd12: n_loc_oh_reg[130] = {3'd0, dist_reg[125], 12'd0};
		4'd13: n_loc_oh_reg[130] = {2'd0, dist_reg[125], 13'd0};
		4'd14: n_loc_oh_reg[130] = {1'd0, dist_reg[125], 14'd0};
		4'd15: n_loc_oh_reg[130] = {dist_reg[125], 15'd0};
	endcase
	case(loc_reg[131])
		4'd0: n_loc_oh_reg[131] = {15'd0, dist_reg[124]};
		4'd1: n_loc_oh_reg[131] = {14'd0, dist_reg[124], 1'd0};
		4'd2: n_loc_oh_reg[131] = {13'd0, dist_reg[124], 2'd0};
		4'd3: n_loc_oh_reg[131] = {12'd0, dist_reg[124], 3'd0};
		4'd4: n_loc_oh_reg[131] = {11'd0, dist_reg[124], 4'd0};
		4'd5: n_loc_oh_reg[131] = {10'd0, dist_reg[124], 5'd0};
		4'd6: n_loc_oh_reg[131] = {9'd0, dist_reg[124], 6'd0};
		4'd7: n_loc_oh_reg[131] = {8'd0, dist_reg[124], 7'd0};
		4'd8: n_loc_oh_reg[131] = {7'd0, dist_reg[124], 8'd0};
		4'd9: n_loc_oh_reg[131] = {6'd0, dist_reg[124], 9'd0};
		4'd10: n_loc_oh_reg[131] = {5'd0, dist_reg[124], 10'd0};
		4'd11: n_loc_oh_reg[131] = {4'd0, dist_reg[124], 11'd0};
		4'd12: n_loc_oh_reg[131] = {3'd0, dist_reg[124], 12'd0};
		4'd13: n_loc_oh_reg[131] = {2'd0, dist_reg[124], 13'd0};
		4'd14: n_loc_oh_reg[131] = {1'd0, dist_reg[124], 14'd0};
		4'd15: n_loc_oh_reg[131] = {dist_reg[124], 15'd0};
	endcase
	case(loc_reg[132])
		4'd0: n_loc_oh_reg[132] = {15'd0, dist_reg[123]};
		4'd1: n_loc_oh_reg[132] = {14'd0, dist_reg[123], 1'd0};
		4'd2: n_loc_oh_reg[132] = {13'd0, dist_reg[123], 2'd0};
		4'd3: n_loc_oh_reg[132] = {12'd0, dist_reg[123], 3'd0};
		4'd4: n_loc_oh_reg[132] = {11'd0, dist_reg[123], 4'd0};
		4'd5: n_loc_oh_reg[132] = {10'd0, dist_reg[123], 5'd0};
		4'd6: n_loc_oh_reg[132] = {9'd0, dist_reg[123], 6'd0};
		4'd7: n_loc_oh_reg[132] = {8'd0, dist_reg[123], 7'd0};
		4'd8: n_loc_oh_reg[132] = {7'd0, dist_reg[123], 8'd0};
		4'd9: n_loc_oh_reg[132] = {6'd0, dist_reg[123], 9'd0};
		4'd10: n_loc_oh_reg[132] = {5'd0, dist_reg[123], 10'd0};
		4'd11: n_loc_oh_reg[132] = {4'd0, dist_reg[123], 11'd0};
		4'd12: n_loc_oh_reg[132] = {3'd0, dist_reg[123], 12'd0};
		4'd13: n_loc_oh_reg[132] = {2'd0, dist_reg[123], 13'd0};
		4'd14: n_loc_oh_reg[132] = {1'd0, dist_reg[123], 14'd0};
		4'd15: n_loc_oh_reg[132] = {dist_reg[123], 15'd0};
	endcase
	case(loc_reg[133])
		4'd0: n_loc_oh_reg[133] = {15'd0, dist_reg[122]};
		4'd1: n_loc_oh_reg[133] = {14'd0, dist_reg[122], 1'd0};
		4'd2: n_loc_oh_reg[133] = {13'd0, dist_reg[122], 2'd0};
		4'd3: n_loc_oh_reg[133] = {12'd0, dist_reg[122], 3'd0};
		4'd4: n_loc_oh_reg[133] = {11'd0, dist_reg[122], 4'd0};
		4'd5: n_loc_oh_reg[133] = {10'd0, dist_reg[122], 5'd0};
		4'd6: n_loc_oh_reg[133] = {9'd0, dist_reg[122], 6'd0};
		4'd7: n_loc_oh_reg[133] = {8'd0, dist_reg[122], 7'd0};
		4'd8: n_loc_oh_reg[133] = {7'd0, dist_reg[122], 8'd0};
		4'd9: n_loc_oh_reg[133] = {6'd0, dist_reg[122], 9'd0};
		4'd10: n_loc_oh_reg[133] = {5'd0, dist_reg[122], 10'd0};
		4'd11: n_loc_oh_reg[133] = {4'd0, dist_reg[122], 11'd0};
		4'd12: n_loc_oh_reg[133] = {3'd0, dist_reg[122], 12'd0};
		4'd13: n_loc_oh_reg[133] = {2'd0, dist_reg[122], 13'd0};
		4'd14: n_loc_oh_reg[133] = {1'd0, dist_reg[122], 14'd0};
		4'd15: n_loc_oh_reg[133] = {dist_reg[122], 15'd0};
	endcase
	case(loc_reg[134])
		4'd0: n_loc_oh_reg[134] = {15'd0, dist_reg[121]};
		4'd1: n_loc_oh_reg[134] = {14'd0, dist_reg[121], 1'd0};
		4'd2: n_loc_oh_reg[134] = {13'd0, dist_reg[121], 2'd0};
		4'd3: n_loc_oh_reg[134] = {12'd0, dist_reg[121], 3'd0};
		4'd4: n_loc_oh_reg[134] = {11'd0, dist_reg[121], 4'd0};
		4'd5: n_loc_oh_reg[134] = {10'd0, dist_reg[121], 5'd0};
		4'd6: n_loc_oh_reg[134] = {9'd0, dist_reg[121], 6'd0};
		4'd7: n_loc_oh_reg[134] = {8'd0, dist_reg[121], 7'd0};
		4'd8: n_loc_oh_reg[134] = {7'd0, dist_reg[121], 8'd0};
		4'd9: n_loc_oh_reg[134] = {6'd0, dist_reg[121], 9'd0};
		4'd10: n_loc_oh_reg[134] = {5'd0, dist_reg[121], 10'd0};
		4'd11: n_loc_oh_reg[134] = {4'd0, dist_reg[121], 11'd0};
		4'd12: n_loc_oh_reg[134] = {3'd0, dist_reg[121], 12'd0};
		4'd13: n_loc_oh_reg[134] = {2'd0, dist_reg[121], 13'd0};
		4'd14: n_loc_oh_reg[134] = {1'd0, dist_reg[121], 14'd0};
		4'd15: n_loc_oh_reg[134] = {dist_reg[121], 15'd0};
	endcase
	case(loc_reg[135])
		4'd0: n_loc_oh_reg[135] = {15'd0, dist_reg[120]};
		4'd1: n_loc_oh_reg[135] = {14'd0, dist_reg[120], 1'd0};
		4'd2: n_loc_oh_reg[135] = {13'd0, dist_reg[120], 2'd0};
		4'd3: n_loc_oh_reg[135] = {12'd0, dist_reg[120], 3'd0};
		4'd4: n_loc_oh_reg[135] = {11'd0, dist_reg[120], 4'd0};
		4'd5: n_loc_oh_reg[135] = {10'd0, dist_reg[120], 5'd0};
		4'd6: n_loc_oh_reg[135] = {9'd0, dist_reg[120], 6'd0};
		4'd7: n_loc_oh_reg[135] = {8'd0, dist_reg[120], 7'd0};
		4'd8: n_loc_oh_reg[135] = {7'd0, dist_reg[120], 8'd0};
		4'd9: n_loc_oh_reg[135] = {6'd0, dist_reg[120], 9'd0};
		4'd10: n_loc_oh_reg[135] = {5'd0, dist_reg[120], 10'd0};
		4'd11: n_loc_oh_reg[135] = {4'd0, dist_reg[120], 11'd0};
		4'd12: n_loc_oh_reg[135] = {3'd0, dist_reg[120], 12'd0};
		4'd13: n_loc_oh_reg[135] = {2'd0, dist_reg[120], 13'd0};
		4'd14: n_loc_oh_reg[135] = {1'd0, dist_reg[120], 14'd0};
		4'd15: n_loc_oh_reg[135] = {dist_reg[120], 15'd0};
	endcase
	case(loc_reg[136])
		4'd0: n_loc_oh_reg[136] = {15'd0, dist_reg[119]};
		4'd1: n_loc_oh_reg[136] = {14'd0, dist_reg[119], 1'd0};
		4'd2: n_loc_oh_reg[136] = {13'd0, dist_reg[119], 2'd0};
		4'd3: n_loc_oh_reg[136] = {12'd0, dist_reg[119], 3'd0};
		4'd4: n_loc_oh_reg[136] = {11'd0, dist_reg[119], 4'd0};
		4'd5: n_loc_oh_reg[136] = {10'd0, dist_reg[119], 5'd0};
		4'd6: n_loc_oh_reg[136] = {9'd0, dist_reg[119], 6'd0};
		4'd7: n_loc_oh_reg[136] = {8'd0, dist_reg[119], 7'd0};
		4'd8: n_loc_oh_reg[136] = {7'd0, dist_reg[119], 8'd0};
		4'd9: n_loc_oh_reg[136] = {6'd0, dist_reg[119], 9'd0};
		4'd10: n_loc_oh_reg[136] = {5'd0, dist_reg[119], 10'd0};
		4'd11: n_loc_oh_reg[136] = {4'd0, dist_reg[119], 11'd0};
		4'd12: n_loc_oh_reg[136] = {3'd0, dist_reg[119], 12'd0};
		4'd13: n_loc_oh_reg[136] = {2'd0, dist_reg[119], 13'd0};
		4'd14: n_loc_oh_reg[136] = {1'd0, dist_reg[119], 14'd0};
		4'd15: n_loc_oh_reg[136] = {dist_reg[119], 15'd0};
	endcase
	case(loc_reg[137])
		4'd0: n_loc_oh_reg[137] = {15'd0, dist_reg[118]};
		4'd1: n_loc_oh_reg[137] = {14'd0, dist_reg[118], 1'd0};
		4'd2: n_loc_oh_reg[137] = {13'd0, dist_reg[118], 2'd0};
		4'd3: n_loc_oh_reg[137] = {12'd0, dist_reg[118], 3'd0};
		4'd4: n_loc_oh_reg[137] = {11'd0, dist_reg[118], 4'd0};
		4'd5: n_loc_oh_reg[137] = {10'd0, dist_reg[118], 5'd0};
		4'd6: n_loc_oh_reg[137] = {9'd0, dist_reg[118], 6'd0};
		4'd7: n_loc_oh_reg[137] = {8'd0, dist_reg[118], 7'd0};
		4'd8: n_loc_oh_reg[137] = {7'd0, dist_reg[118], 8'd0};
		4'd9: n_loc_oh_reg[137] = {6'd0, dist_reg[118], 9'd0};
		4'd10: n_loc_oh_reg[137] = {5'd0, dist_reg[118], 10'd0};
		4'd11: n_loc_oh_reg[137] = {4'd0, dist_reg[118], 11'd0};
		4'd12: n_loc_oh_reg[137] = {3'd0, dist_reg[118], 12'd0};
		4'd13: n_loc_oh_reg[137] = {2'd0, dist_reg[118], 13'd0};
		4'd14: n_loc_oh_reg[137] = {1'd0, dist_reg[118], 14'd0};
		4'd15: n_loc_oh_reg[137] = {dist_reg[118], 15'd0};
	endcase
	case(loc_reg[138])
		4'd0: n_loc_oh_reg[138] = {15'd0, dist_reg[117]};
		4'd1: n_loc_oh_reg[138] = {14'd0, dist_reg[117], 1'd0};
		4'd2: n_loc_oh_reg[138] = {13'd0, dist_reg[117], 2'd0};
		4'd3: n_loc_oh_reg[138] = {12'd0, dist_reg[117], 3'd0};
		4'd4: n_loc_oh_reg[138] = {11'd0, dist_reg[117], 4'd0};
		4'd5: n_loc_oh_reg[138] = {10'd0, dist_reg[117], 5'd0};
		4'd6: n_loc_oh_reg[138] = {9'd0, dist_reg[117], 6'd0};
		4'd7: n_loc_oh_reg[138] = {8'd0, dist_reg[117], 7'd0};
		4'd8: n_loc_oh_reg[138] = {7'd0, dist_reg[117], 8'd0};
		4'd9: n_loc_oh_reg[138] = {6'd0, dist_reg[117], 9'd0};
		4'd10: n_loc_oh_reg[138] = {5'd0, dist_reg[117], 10'd0};
		4'd11: n_loc_oh_reg[138] = {4'd0, dist_reg[117], 11'd0};
		4'd12: n_loc_oh_reg[138] = {3'd0, dist_reg[117], 12'd0};
		4'd13: n_loc_oh_reg[138] = {2'd0, dist_reg[117], 13'd0};
		4'd14: n_loc_oh_reg[138] = {1'd0, dist_reg[117], 14'd0};
		4'd15: n_loc_oh_reg[138] = {dist_reg[117], 15'd0};
	endcase
	case(loc_reg[139])
		4'd0: n_loc_oh_reg[139] = {15'd0, dist_reg[116]};
		4'd1: n_loc_oh_reg[139] = {14'd0, dist_reg[116], 1'd0};
		4'd2: n_loc_oh_reg[139] = {13'd0, dist_reg[116], 2'd0};
		4'd3: n_loc_oh_reg[139] = {12'd0, dist_reg[116], 3'd0};
		4'd4: n_loc_oh_reg[139] = {11'd0, dist_reg[116], 4'd0};
		4'd5: n_loc_oh_reg[139] = {10'd0, dist_reg[116], 5'd0};
		4'd6: n_loc_oh_reg[139] = {9'd0, dist_reg[116], 6'd0};
		4'd7: n_loc_oh_reg[139] = {8'd0, dist_reg[116], 7'd0};
		4'd8: n_loc_oh_reg[139] = {7'd0, dist_reg[116], 8'd0};
		4'd9: n_loc_oh_reg[139] = {6'd0, dist_reg[116], 9'd0};
		4'd10: n_loc_oh_reg[139] = {5'd0, dist_reg[116], 10'd0};
		4'd11: n_loc_oh_reg[139] = {4'd0, dist_reg[116], 11'd0};
		4'd12: n_loc_oh_reg[139] = {3'd0, dist_reg[116], 12'd0};
		4'd13: n_loc_oh_reg[139] = {2'd0, dist_reg[116], 13'd0};
		4'd14: n_loc_oh_reg[139] = {1'd0, dist_reg[116], 14'd0};
		4'd15: n_loc_oh_reg[139] = {dist_reg[116], 15'd0};
	endcase
	case(loc_reg[140])
		4'd0: n_loc_oh_reg[140] = {15'd0, dist_reg[115]};
		4'd1: n_loc_oh_reg[140] = {14'd0, dist_reg[115], 1'd0};
		4'd2: n_loc_oh_reg[140] = {13'd0, dist_reg[115], 2'd0};
		4'd3: n_loc_oh_reg[140] = {12'd0, dist_reg[115], 3'd0};
		4'd4: n_loc_oh_reg[140] = {11'd0, dist_reg[115], 4'd0};
		4'd5: n_loc_oh_reg[140] = {10'd0, dist_reg[115], 5'd0};
		4'd6: n_loc_oh_reg[140] = {9'd0, dist_reg[115], 6'd0};
		4'd7: n_loc_oh_reg[140] = {8'd0, dist_reg[115], 7'd0};
		4'd8: n_loc_oh_reg[140] = {7'd0, dist_reg[115], 8'd0};
		4'd9: n_loc_oh_reg[140] = {6'd0, dist_reg[115], 9'd0};
		4'd10: n_loc_oh_reg[140] = {5'd0, dist_reg[115], 10'd0};
		4'd11: n_loc_oh_reg[140] = {4'd0, dist_reg[115], 11'd0};
		4'd12: n_loc_oh_reg[140] = {3'd0, dist_reg[115], 12'd0};
		4'd13: n_loc_oh_reg[140] = {2'd0, dist_reg[115], 13'd0};
		4'd14: n_loc_oh_reg[140] = {1'd0, dist_reg[115], 14'd0};
		4'd15: n_loc_oh_reg[140] = {dist_reg[115], 15'd0};
	endcase
	case(loc_reg[141])
		4'd0: n_loc_oh_reg[141] = {15'd0, dist_reg[114]};
		4'd1: n_loc_oh_reg[141] = {14'd0, dist_reg[114], 1'd0};
		4'd2: n_loc_oh_reg[141] = {13'd0, dist_reg[114], 2'd0};
		4'd3: n_loc_oh_reg[141] = {12'd0, dist_reg[114], 3'd0};
		4'd4: n_loc_oh_reg[141] = {11'd0, dist_reg[114], 4'd0};
		4'd5: n_loc_oh_reg[141] = {10'd0, dist_reg[114], 5'd0};
		4'd6: n_loc_oh_reg[141] = {9'd0, dist_reg[114], 6'd0};
		4'd7: n_loc_oh_reg[141] = {8'd0, dist_reg[114], 7'd0};
		4'd8: n_loc_oh_reg[141] = {7'd0, dist_reg[114], 8'd0};
		4'd9: n_loc_oh_reg[141] = {6'd0, dist_reg[114], 9'd0};
		4'd10: n_loc_oh_reg[141] = {5'd0, dist_reg[114], 10'd0};
		4'd11: n_loc_oh_reg[141] = {4'd0, dist_reg[114], 11'd0};
		4'd12: n_loc_oh_reg[141] = {3'd0, dist_reg[114], 12'd0};
		4'd13: n_loc_oh_reg[141] = {2'd0, dist_reg[114], 13'd0};
		4'd14: n_loc_oh_reg[141] = {1'd0, dist_reg[114], 14'd0};
		4'd15: n_loc_oh_reg[141] = {dist_reg[114], 15'd0};
	endcase
	case(loc_reg[142])
		4'd0: n_loc_oh_reg[142] = {15'd0, dist_reg[113]};
		4'd1: n_loc_oh_reg[142] = {14'd0, dist_reg[113], 1'd0};
		4'd2: n_loc_oh_reg[142] = {13'd0, dist_reg[113], 2'd0};
		4'd3: n_loc_oh_reg[142] = {12'd0, dist_reg[113], 3'd0};
		4'd4: n_loc_oh_reg[142] = {11'd0, dist_reg[113], 4'd0};
		4'd5: n_loc_oh_reg[142] = {10'd0, dist_reg[113], 5'd0};
		4'd6: n_loc_oh_reg[142] = {9'd0, dist_reg[113], 6'd0};
		4'd7: n_loc_oh_reg[142] = {8'd0, dist_reg[113], 7'd0};
		4'd8: n_loc_oh_reg[142] = {7'd0, dist_reg[113], 8'd0};
		4'd9: n_loc_oh_reg[142] = {6'd0, dist_reg[113], 9'd0};
		4'd10: n_loc_oh_reg[142] = {5'd0, dist_reg[113], 10'd0};
		4'd11: n_loc_oh_reg[142] = {4'd0, dist_reg[113], 11'd0};
		4'd12: n_loc_oh_reg[142] = {3'd0, dist_reg[113], 12'd0};
		4'd13: n_loc_oh_reg[142] = {2'd0, dist_reg[113], 13'd0};
		4'd14: n_loc_oh_reg[142] = {1'd0, dist_reg[113], 14'd0};
		4'd15: n_loc_oh_reg[142] = {dist_reg[113], 15'd0};
	endcase
	case(loc_reg[143])
		4'd0: n_loc_oh_reg[143] = {15'd0, dist_reg[112]};
		4'd1: n_loc_oh_reg[143] = {14'd0, dist_reg[112], 1'd0};
		4'd2: n_loc_oh_reg[143] = {13'd0, dist_reg[112], 2'd0};
		4'd3: n_loc_oh_reg[143] = {12'd0, dist_reg[112], 3'd0};
		4'd4: n_loc_oh_reg[143] = {11'd0, dist_reg[112], 4'd0};
		4'd5: n_loc_oh_reg[143] = {10'd0, dist_reg[112], 5'd0};
		4'd6: n_loc_oh_reg[143] = {9'd0, dist_reg[112], 6'd0};
		4'd7: n_loc_oh_reg[143] = {8'd0, dist_reg[112], 7'd0};
		4'd8: n_loc_oh_reg[143] = {7'd0, dist_reg[112], 8'd0};
		4'd9: n_loc_oh_reg[143] = {6'd0, dist_reg[112], 9'd0};
		4'd10: n_loc_oh_reg[143] = {5'd0, dist_reg[112], 10'd0};
		4'd11: n_loc_oh_reg[143] = {4'd0, dist_reg[112], 11'd0};
		4'd12: n_loc_oh_reg[143] = {3'd0, dist_reg[112], 12'd0};
		4'd13: n_loc_oh_reg[143] = {2'd0, dist_reg[112], 13'd0};
		4'd14: n_loc_oh_reg[143] = {1'd0, dist_reg[112], 14'd0};
		4'd15: n_loc_oh_reg[143] = {dist_reg[112], 15'd0};
	endcase
	case(loc_reg[144])
		4'd0: n_loc_oh_reg[144] = {15'd0, dist_reg[111]};
		4'd1: n_loc_oh_reg[144] = {14'd0, dist_reg[111], 1'd0};
		4'd2: n_loc_oh_reg[144] = {13'd0, dist_reg[111], 2'd0};
		4'd3: n_loc_oh_reg[144] = {12'd0, dist_reg[111], 3'd0};
		4'd4: n_loc_oh_reg[144] = {11'd0, dist_reg[111], 4'd0};
		4'd5: n_loc_oh_reg[144] = {10'd0, dist_reg[111], 5'd0};
		4'd6: n_loc_oh_reg[144] = {9'd0, dist_reg[111], 6'd0};
		4'd7: n_loc_oh_reg[144] = {8'd0, dist_reg[111], 7'd0};
		4'd8: n_loc_oh_reg[144] = {7'd0, dist_reg[111], 8'd0};
		4'd9: n_loc_oh_reg[144] = {6'd0, dist_reg[111], 9'd0};
		4'd10: n_loc_oh_reg[144] = {5'd0, dist_reg[111], 10'd0};
		4'd11: n_loc_oh_reg[144] = {4'd0, dist_reg[111], 11'd0};
		4'd12: n_loc_oh_reg[144] = {3'd0, dist_reg[111], 12'd0};
		4'd13: n_loc_oh_reg[144] = {2'd0, dist_reg[111], 13'd0};
		4'd14: n_loc_oh_reg[144] = {1'd0, dist_reg[111], 14'd0};
		4'd15: n_loc_oh_reg[144] = {dist_reg[111], 15'd0};
	endcase
	case(loc_reg[145])
		4'd0: n_loc_oh_reg[145] = {15'd0, dist_reg[110]};
		4'd1: n_loc_oh_reg[145] = {14'd0, dist_reg[110], 1'd0};
		4'd2: n_loc_oh_reg[145] = {13'd0, dist_reg[110], 2'd0};
		4'd3: n_loc_oh_reg[145] = {12'd0, dist_reg[110], 3'd0};
		4'd4: n_loc_oh_reg[145] = {11'd0, dist_reg[110], 4'd0};
		4'd5: n_loc_oh_reg[145] = {10'd0, dist_reg[110], 5'd0};
		4'd6: n_loc_oh_reg[145] = {9'd0, dist_reg[110], 6'd0};
		4'd7: n_loc_oh_reg[145] = {8'd0, dist_reg[110], 7'd0};
		4'd8: n_loc_oh_reg[145] = {7'd0, dist_reg[110], 8'd0};
		4'd9: n_loc_oh_reg[145] = {6'd0, dist_reg[110], 9'd0};
		4'd10: n_loc_oh_reg[145] = {5'd0, dist_reg[110], 10'd0};
		4'd11: n_loc_oh_reg[145] = {4'd0, dist_reg[110], 11'd0};
		4'd12: n_loc_oh_reg[145] = {3'd0, dist_reg[110], 12'd0};
		4'd13: n_loc_oh_reg[145] = {2'd0, dist_reg[110], 13'd0};
		4'd14: n_loc_oh_reg[145] = {1'd0, dist_reg[110], 14'd0};
		4'd15: n_loc_oh_reg[145] = {dist_reg[110], 15'd0};
	endcase
	case(loc_reg[146])
		4'd0: n_loc_oh_reg[146] = {15'd0, dist_reg[109]};
		4'd1: n_loc_oh_reg[146] = {14'd0, dist_reg[109], 1'd0};
		4'd2: n_loc_oh_reg[146] = {13'd0, dist_reg[109], 2'd0};
		4'd3: n_loc_oh_reg[146] = {12'd0, dist_reg[109], 3'd0};
		4'd4: n_loc_oh_reg[146] = {11'd0, dist_reg[109], 4'd0};
		4'd5: n_loc_oh_reg[146] = {10'd0, dist_reg[109], 5'd0};
		4'd6: n_loc_oh_reg[146] = {9'd0, dist_reg[109], 6'd0};
		4'd7: n_loc_oh_reg[146] = {8'd0, dist_reg[109], 7'd0};
		4'd8: n_loc_oh_reg[146] = {7'd0, dist_reg[109], 8'd0};
		4'd9: n_loc_oh_reg[146] = {6'd0, dist_reg[109], 9'd0};
		4'd10: n_loc_oh_reg[146] = {5'd0, dist_reg[109], 10'd0};
		4'd11: n_loc_oh_reg[146] = {4'd0, dist_reg[109], 11'd0};
		4'd12: n_loc_oh_reg[146] = {3'd0, dist_reg[109], 12'd0};
		4'd13: n_loc_oh_reg[146] = {2'd0, dist_reg[109], 13'd0};
		4'd14: n_loc_oh_reg[146] = {1'd0, dist_reg[109], 14'd0};
		4'd15: n_loc_oh_reg[146] = {dist_reg[109], 15'd0};
	endcase
	case(loc_reg[147])
		4'd0: n_loc_oh_reg[147] = {15'd0, dist_reg[108]};
		4'd1: n_loc_oh_reg[147] = {14'd0, dist_reg[108], 1'd0};
		4'd2: n_loc_oh_reg[147] = {13'd0, dist_reg[108], 2'd0};
		4'd3: n_loc_oh_reg[147] = {12'd0, dist_reg[108], 3'd0};
		4'd4: n_loc_oh_reg[147] = {11'd0, dist_reg[108], 4'd0};
		4'd5: n_loc_oh_reg[147] = {10'd0, dist_reg[108], 5'd0};
		4'd6: n_loc_oh_reg[147] = {9'd0, dist_reg[108], 6'd0};
		4'd7: n_loc_oh_reg[147] = {8'd0, dist_reg[108], 7'd0};
		4'd8: n_loc_oh_reg[147] = {7'd0, dist_reg[108], 8'd0};
		4'd9: n_loc_oh_reg[147] = {6'd0, dist_reg[108], 9'd0};
		4'd10: n_loc_oh_reg[147] = {5'd0, dist_reg[108], 10'd0};
		4'd11: n_loc_oh_reg[147] = {4'd0, dist_reg[108], 11'd0};
		4'd12: n_loc_oh_reg[147] = {3'd0, dist_reg[108], 12'd0};
		4'd13: n_loc_oh_reg[147] = {2'd0, dist_reg[108], 13'd0};
		4'd14: n_loc_oh_reg[147] = {1'd0, dist_reg[108], 14'd0};
		4'd15: n_loc_oh_reg[147] = {dist_reg[108], 15'd0};
	endcase
	case(loc_reg[148])
		4'd0: n_loc_oh_reg[148] = {15'd0, dist_reg[107]};
		4'd1: n_loc_oh_reg[148] = {14'd0, dist_reg[107], 1'd0};
		4'd2: n_loc_oh_reg[148] = {13'd0, dist_reg[107], 2'd0};
		4'd3: n_loc_oh_reg[148] = {12'd0, dist_reg[107], 3'd0};
		4'd4: n_loc_oh_reg[148] = {11'd0, dist_reg[107], 4'd0};
		4'd5: n_loc_oh_reg[148] = {10'd0, dist_reg[107], 5'd0};
		4'd6: n_loc_oh_reg[148] = {9'd0, dist_reg[107], 6'd0};
		4'd7: n_loc_oh_reg[148] = {8'd0, dist_reg[107], 7'd0};
		4'd8: n_loc_oh_reg[148] = {7'd0, dist_reg[107], 8'd0};
		4'd9: n_loc_oh_reg[148] = {6'd0, dist_reg[107], 9'd0};
		4'd10: n_loc_oh_reg[148] = {5'd0, dist_reg[107], 10'd0};
		4'd11: n_loc_oh_reg[148] = {4'd0, dist_reg[107], 11'd0};
		4'd12: n_loc_oh_reg[148] = {3'd0, dist_reg[107], 12'd0};
		4'd13: n_loc_oh_reg[148] = {2'd0, dist_reg[107], 13'd0};
		4'd14: n_loc_oh_reg[148] = {1'd0, dist_reg[107], 14'd0};
		4'd15: n_loc_oh_reg[148] = {dist_reg[107], 15'd0};
	endcase
	case(loc_reg[149])
		4'd0: n_loc_oh_reg[149] = {15'd0, dist_reg[106]};
		4'd1: n_loc_oh_reg[149] = {14'd0, dist_reg[106], 1'd0};
		4'd2: n_loc_oh_reg[149] = {13'd0, dist_reg[106], 2'd0};
		4'd3: n_loc_oh_reg[149] = {12'd0, dist_reg[106], 3'd0};
		4'd4: n_loc_oh_reg[149] = {11'd0, dist_reg[106], 4'd0};
		4'd5: n_loc_oh_reg[149] = {10'd0, dist_reg[106], 5'd0};
		4'd6: n_loc_oh_reg[149] = {9'd0, dist_reg[106], 6'd0};
		4'd7: n_loc_oh_reg[149] = {8'd0, dist_reg[106], 7'd0};
		4'd8: n_loc_oh_reg[149] = {7'd0, dist_reg[106], 8'd0};
		4'd9: n_loc_oh_reg[149] = {6'd0, dist_reg[106], 9'd0};
		4'd10: n_loc_oh_reg[149] = {5'd0, dist_reg[106], 10'd0};
		4'd11: n_loc_oh_reg[149] = {4'd0, dist_reg[106], 11'd0};
		4'd12: n_loc_oh_reg[149] = {3'd0, dist_reg[106], 12'd0};
		4'd13: n_loc_oh_reg[149] = {2'd0, dist_reg[106], 13'd0};
		4'd14: n_loc_oh_reg[149] = {1'd0, dist_reg[106], 14'd0};
		4'd15: n_loc_oh_reg[149] = {dist_reg[106], 15'd0};
	endcase
	case(loc_reg[150])
		4'd0: n_loc_oh_reg[150] = {15'd0, dist_reg[105]};
		4'd1: n_loc_oh_reg[150] = {14'd0, dist_reg[105], 1'd0};
		4'd2: n_loc_oh_reg[150] = {13'd0, dist_reg[105], 2'd0};
		4'd3: n_loc_oh_reg[150] = {12'd0, dist_reg[105], 3'd0};
		4'd4: n_loc_oh_reg[150] = {11'd0, dist_reg[105], 4'd0};
		4'd5: n_loc_oh_reg[150] = {10'd0, dist_reg[105], 5'd0};
		4'd6: n_loc_oh_reg[150] = {9'd0, dist_reg[105], 6'd0};
		4'd7: n_loc_oh_reg[150] = {8'd0, dist_reg[105], 7'd0};
		4'd8: n_loc_oh_reg[150] = {7'd0, dist_reg[105], 8'd0};
		4'd9: n_loc_oh_reg[150] = {6'd0, dist_reg[105], 9'd0};
		4'd10: n_loc_oh_reg[150] = {5'd0, dist_reg[105], 10'd0};
		4'd11: n_loc_oh_reg[150] = {4'd0, dist_reg[105], 11'd0};
		4'd12: n_loc_oh_reg[150] = {3'd0, dist_reg[105], 12'd0};
		4'd13: n_loc_oh_reg[150] = {2'd0, dist_reg[105], 13'd0};
		4'd14: n_loc_oh_reg[150] = {1'd0, dist_reg[105], 14'd0};
		4'd15: n_loc_oh_reg[150] = {dist_reg[105], 15'd0};
	endcase
	case(loc_reg[151])
		4'd0: n_loc_oh_reg[151] = {15'd0, dist_reg[104]};
		4'd1: n_loc_oh_reg[151] = {14'd0, dist_reg[104], 1'd0};
		4'd2: n_loc_oh_reg[151] = {13'd0, dist_reg[104], 2'd0};
		4'd3: n_loc_oh_reg[151] = {12'd0, dist_reg[104], 3'd0};
		4'd4: n_loc_oh_reg[151] = {11'd0, dist_reg[104], 4'd0};
		4'd5: n_loc_oh_reg[151] = {10'd0, dist_reg[104], 5'd0};
		4'd6: n_loc_oh_reg[151] = {9'd0, dist_reg[104], 6'd0};
		4'd7: n_loc_oh_reg[151] = {8'd0, dist_reg[104], 7'd0};
		4'd8: n_loc_oh_reg[151] = {7'd0, dist_reg[104], 8'd0};
		4'd9: n_loc_oh_reg[151] = {6'd0, dist_reg[104], 9'd0};
		4'd10: n_loc_oh_reg[151] = {5'd0, dist_reg[104], 10'd0};
		4'd11: n_loc_oh_reg[151] = {4'd0, dist_reg[104], 11'd0};
		4'd12: n_loc_oh_reg[151] = {3'd0, dist_reg[104], 12'd0};
		4'd13: n_loc_oh_reg[151] = {2'd0, dist_reg[104], 13'd0};
		4'd14: n_loc_oh_reg[151] = {1'd0, dist_reg[104], 14'd0};
		4'd15: n_loc_oh_reg[151] = {dist_reg[104], 15'd0};
	endcase
	case(loc_reg[152])
		4'd0: n_loc_oh_reg[152] = {15'd0, dist_reg[103]};
		4'd1: n_loc_oh_reg[152] = {14'd0, dist_reg[103], 1'd0};
		4'd2: n_loc_oh_reg[152] = {13'd0, dist_reg[103], 2'd0};
		4'd3: n_loc_oh_reg[152] = {12'd0, dist_reg[103], 3'd0};
		4'd4: n_loc_oh_reg[152] = {11'd0, dist_reg[103], 4'd0};
		4'd5: n_loc_oh_reg[152] = {10'd0, dist_reg[103], 5'd0};
		4'd6: n_loc_oh_reg[152] = {9'd0, dist_reg[103], 6'd0};
		4'd7: n_loc_oh_reg[152] = {8'd0, dist_reg[103], 7'd0};
		4'd8: n_loc_oh_reg[152] = {7'd0, dist_reg[103], 8'd0};
		4'd9: n_loc_oh_reg[152] = {6'd0, dist_reg[103], 9'd0};
		4'd10: n_loc_oh_reg[152] = {5'd0, dist_reg[103], 10'd0};
		4'd11: n_loc_oh_reg[152] = {4'd0, dist_reg[103], 11'd0};
		4'd12: n_loc_oh_reg[152] = {3'd0, dist_reg[103], 12'd0};
		4'd13: n_loc_oh_reg[152] = {2'd0, dist_reg[103], 13'd0};
		4'd14: n_loc_oh_reg[152] = {1'd0, dist_reg[103], 14'd0};
		4'd15: n_loc_oh_reg[152] = {dist_reg[103], 15'd0};
	endcase
	case(loc_reg[153])
		4'd0: n_loc_oh_reg[153] = {15'd0, dist_reg[102]};
		4'd1: n_loc_oh_reg[153] = {14'd0, dist_reg[102], 1'd0};
		4'd2: n_loc_oh_reg[153] = {13'd0, dist_reg[102], 2'd0};
		4'd3: n_loc_oh_reg[153] = {12'd0, dist_reg[102], 3'd0};
		4'd4: n_loc_oh_reg[153] = {11'd0, dist_reg[102], 4'd0};
		4'd5: n_loc_oh_reg[153] = {10'd0, dist_reg[102], 5'd0};
		4'd6: n_loc_oh_reg[153] = {9'd0, dist_reg[102], 6'd0};
		4'd7: n_loc_oh_reg[153] = {8'd0, dist_reg[102], 7'd0};
		4'd8: n_loc_oh_reg[153] = {7'd0, dist_reg[102], 8'd0};
		4'd9: n_loc_oh_reg[153] = {6'd0, dist_reg[102], 9'd0};
		4'd10: n_loc_oh_reg[153] = {5'd0, dist_reg[102], 10'd0};
		4'd11: n_loc_oh_reg[153] = {4'd0, dist_reg[102], 11'd0};
		4'd12: n_loc_oh_reg[153] = {3'd0, dist_reg[102], 12'd0};
		4'd13: n_loc_oh_reg[153] = {2'd0, dist_reg[102], 13'd0};
		4'd14: n_loc_oh_reg[153] = {1'd0, dist_reg[102], 14'd0};
		4'd15: n_loc_oh_reg[153] = {dist_reg[102], 15'd0};
	endcase
	case(loc_reg[154])
		4'd0: n_loc_oh_reg[154] = {15'd0, dist_reg[101]};
		4'd1: n_loc_oh_reg[154] = {14'd0, dist_reg[101], 1'd0};
		4'd2: n_loc_oh_reg[154] = {13'd0, dist_reg[101], 2'd0};
		4'd3: n_loc_oh_reg[154] = {12'd0, dist_reg[101], 3'd0};
		4'd4: n_loc_oh_reg[154] = {11'd0, dist_reg[101], 4'd0};
		4'd5: n_loc_oh_reg[154] = {10'd0, dist_reg[101], 5'd0};
		4'd6: n_loc_oh_reg[154] = {9'd0, dist_reg[101], 6'd0};
		4'd7: n_loc_oh_reg[154] = {8'd0, dist_reg[101], 7'd0};
		4'd8: n_loc_oh_reg[154] = {7'd0, dist_reg[101], 8'd0};
		4'd9: n_loc_oh_reg[154] = {6'd0, dist_reg[101], 9'd0};
		4'd10: n_loc_oh_reg[154] = {5'd0, dist_reg[101], 10'd0};
		4'd11: n_loc_oh_reg[154] = {4'd0, dist_reg[101], 11'd0};
		4'd12: n_loc_oh_reg[154] = {3'd0, dist_reg[101], 12'd0};
		4'd13: n_loc_oh_reg[154] = {2'd0, dist_reg[101], 13'd0};
		4'd14: n_loc_oh_reg[154] = {1'd0, dist_reg[101], 14'd0};
		4'd15: n_loc_oh_reg[154] = {dist_reg[101], 15'd0};
	endcase
	case(loc_reg[155])
		4'd0: n_loc_oh_reg[155] = {15'd0, dist_reg[100]};
		4'd1: n_loc_oh_reg[155] = {14'd0, dist_reg[100], 1'd0};
		4'd2: n_loc_oh_reg[155] = {13'd0, dist_reg[100], 2'd0};
		4'd3: n_loc_oh_reg[155] = {12'd0, dist_reg[100], 3'd0};
		4'd4: n_loc_oh_reg[155] = {11'd0, dist_reg[100], 4'd0};
		4'd5: n_loc_oh_reg[155] = {10'd0, dist_reg[100], 5'd0};
		4'd6: n_loc_oh_reg[155] = {9'd0, dist_reg[100], 6'd0};
		4'd7: n_loc_oh_reg[155] = {8'd0, dist_reg[100], 7'd0};
		4'd8: n_loc_oh_reg[155] = {7'd0, dist_reg[100], 8'd0};
		4'd9: n_loc_oh_reg[155] = {6'd0, dist_reg[100], 9'd0};
		4'd10: n_loc_oh_reg[155] = {5'd0, dist_reg[100], 10'd0};
		4'd11: n_loc_oh_reg[155] = {4'd0, dist_reg[100], 11'd0};
		4'd12: n_loc_oh_reg[155] = {3'd0, dist_reg[100], 12'd0};
		4'd13: n_loc_oh_reg[155] = {2'd0, dist_reg[100], 13'd0};
		4'd14: n_loc_oh_reg[155] = {1'd0, dist_reg[100], 14'd0};
		4'd15: n_loc_oh_reg[155] = {dist_reg[100], 15'd0};
	endcase
	case(loc_reg[156])
		4'd0: n_loc_oh_reg[156] = {15'd0, dist_reg[99]};
		4'd1: n_loc_oh_reg[156] = {14'd0, dist_reg[99], 1'd0};
		4'd2: n_loc_oh_reg[156] = {13'd0, dist_reg[99], 2'd0};
		4'd3: n_loc_oh_reg[156] = {12'd0, dist_reg[99], 3'd0};
		4'd4: n_loc_oh_reg[156] = {11'd0, dist_reg[99], 4'd0};
		4'd5: n_loc_oh_reg[156] = {10'd0, dist_reg[99], 5'd0};
		4'd6: n_loc_oh_reg[156] = {9'd0, dist_reg[99], 6'd0};
		4'd7: n_loc_oh_reg[156] = {8'd0, dist_reg[99], 7'd0};
		4'd8: n_loc_oh_reg[156] = {7'd0, dist_reg[99], 8'd0};
		4'd9: n_loc_oh_reg[156] = {6'd0, dist_reg[99], 9'd0};
		4'd10: n_loc_oh_reg[156] = {5'd0, dist_reg[99], 10'd0};
		4'd11: n_loc_oh_reg[156] = {4'd0, dist_reg[99], 11'd0};
		4'd12: n_loc_oh_reg[156] = {3'd0, dist_reg[99], 12'd0};
		4'd13: n_loc_oh_reg[156] = {2'd0, dist_reg[99], 13'd0};
		4'd14: n_loc_oh_reg[156] = {1'd0, dist_reg[99], 14'd0};
		4'd15: n_loc_oh_reg[156] = {dist_reg[99], 15'd0};
	endcase
	case(loc_reg[157])
		4'd0: n_loc_oh_reg[157] = {15'd0, dist_reg[98]};
		4'd1: n_loc_oh_reg[157] = {14'd0, dist_reg[98], 1'd0};
		4'd2: n_loc_oh_reg[157] = {13'd0, dist_reg[98], 2'd0};
		4'd3: n_loc_oh_reg[157] = {12'd0, dist_reg[98], 3'd0};
		4'd4: n_loc_oh_reg[157] = {11'd0, dist_reg[98], 4'd0};
		4'd5: n_loc_oh_reg[157] = {10'd0, dist_reg[98], 5'd0};
		4'd6: n_loc_oh_reg[157] = {9'd0, dist_reg[98], 6'd0};
		4'd7: n_loc_oh_reg[157] = {8'd0, dist_reg[98], 7'd0};
		4'd8: n_loc_oh_reg[157] = {7'd0, dist_reg[98], 8'd0};
		4'd9: n_loc_oh_reg[157] = {6'd0, dist_reg[98], 9'd0};
		4'd10: n_loc_oh_reg[157] = {5'd0, dist_reg[98], 10'd0};
		4'd11: n_loc_oh_reg[157] = {4'd0, dist_reg[98], 11'd0};
		4'd12: n_loc_oh_reg[157] = {3'd0, dist_reg[98], 12'd0};
		4'd13: n_loc_oh_reg[157] = {2'd0, dist_reg[98], 13'd0};
		4'd14: n_loc_oh_reg[157] = {1'd0, dist_reg[98], 14'd0};
		4'd15: n_loc_oh_reg[157] = {dist_reg[98], 15'd0};
	endcase
	case(loc_reg[158])
		4'd0: n_loc_oh_reg[158] = {15'd0, dist_reg[97]};
		4'd1: n_loc_oh_reg[158] = {14'd0, dist_reg[97], 1'd0};
		4'd2: n_loc_oh_reg[158] = {13'd0, dist_reg[97], 2'd0};
		4'd3: n_loc_oh_reg[158] = {12'd0, dist_reg[97], 3'd0};
		4'd4: n_loc_oh_reg[158] = {11'd0, dist_reg[97], 4'd0};
		4'd5: n_loc_oh_reg[158] = {10'd0, dist_reg[97], 5'd0};
		4'd6: n_loc_oh_reg[158] = {9'd0, dist_reg[97], 6'd0};
		4'd7: n_loc_oh_reg[158] = {8'd0, dist_reg[97], 7'd0};
		4'd8: n_loc_oh_reg[158] = {7'd0, dist_reg[97], 8'd0};
		4'd9: n_loc_oh_reg[158] = {6'd0, dist_reg[97], 9'd0};
		4'd10: n_loc_oh_reg[158] = {5'd0, dist_reg[97], 10'd0};
		4'd11: n_loc_oh_reg[158] = {4'd0, dist_reg[97], 11'd0};
		4'd12: n_loc_oh_reg[158] = {3'd0, dist_reg[97], 12'd0};
		4'd13: n_loc_oh_reg[158] = {2'd0, dist_reg[97], 13'd0};
		4'd14: n_loc_oh_reg[158] = {1'd0, dist_reg[97], 14'd0};
		4'd15: n_loc_oh_reg[158] = {dist_reg[97], 15'd0};
	endcase
	case(loc_reg[159])
		4'd0: n_loc_oh_reg[159] = {15'd0, dist_reg[96]};
		4'd1: n_loc_oh_reg[159] = {14'd0, dist_reg[96], 1'd0};
		4'd2: n_loc_oh_reg[159] = {13'd0, dist_reg[96], 2'd0};
		4'd3: n_loc_oh_reg[159] = {12'd0, dist_reg[96], 3'd0};
		4'd4: n_loc_oh_reg[159] = {11'd0, dist_reg[96], 4'd0};
		4'd5: n_loc_oh_reg[159] = {10'd0, dist_reg[96], 5'd0};
		4'd6: n_loc_oh_reg[159] = {9'd0, dist_reg[96], 6'd0};
		4'd7: n_loc_oh_reg[159] = {8'd0, dist_reg[96], 7'd0};
		4'd8: n_loc_oh_reg[159] = {7'd0, dist_reg[96], 8'd0};
		4'd9: n_loc_oh_reg[159] = {6'd0, dist_reg[96], 9'd0};
		4'd10: n_loc_oh_reg[159] = {5'd0, dist_reg[96], 10'd0};
		4'd11: n_loc_oh_reg[159] = {4'd0, dist_reg[96], 11'd0};
		4'd12: n_loc_oh_reg[159] = {3'd0, dist_reg[96], 12'd0};
		4'd13: n_loc_oh_reg[159] = {2'd0, dist_reg[96], 13'd0};
		4'd14: n_loc_oh_reg[159] = {1'd0, dist_reg[96], 14'd0};
		4'd15: n_loc_oh_reg[159] = {dist_reg[96], 15'd0};
	endcase
	case(loc_reg[160])
		4'd0: n_loc_oh_reg[160] = {15'd0, dist_reg[95]};
		4'd1: n_loc_oh_reg[160] = {14'd0, dist_reg[95], 1'd0};
		4'd2: n_loc_oh_reg[160] = {13'd0, dist_reg[95], 2'd0};
		4'd3: n_loc_oh_reg[160] = {12'd0, dist_reg[95], 3'd0};
		4'd4: n_loc_oh_reg[160] = {11'd0, dist_reg[95], 4'd0};
		4'd5: n_loc_oh_reg[160] = {10'd0, dist_reg[95], 5'd0};
		4'd6: n_loc_oh_reg[160] = {9'd0, dist_reg[95], 6'd0};
		4'd7: n_loc_oh_reg[160] = {8'd0, dist_reg[95], 7'd0};
		4'd8: n_loc_oh_reg[160] = {7'd0, dist_reg[95], 8'd0};
		4'd9: n_loc_oh_reg[160] = {6'd0, dist_reg[95], 9'd0};
		4'd10: n_loc_oh_reg[160] = {5'd0, dist_reg[95], 10'd0};
		4'd11: n_loc_oh_reg[160] = {4'd0, dist_reg[95], 11'd0};
		4'd12: n_loc_oh_reg[160] = {3'd0, dist_reg[95], 12'd0};
		4'd13: n_loc_oh_reg[160] = {2'd0, dist_reg[95], 13'd0};
		4'd14: n_loc_oh_reg[160] = {1'd0, dist_reg[95], 14'd0};
		4'd15: n_loc_oh_reg[160] = {dist_reg[95], 15'd0};
	endcase
	case(loc_reg[161])
		4'd0: n_loc_oh_reg[161] = {15'd0, dist_reg[94]};
		4'd1: n_loc_oh_reg[161] = {14'd0, dist_reg[94], 1'd0};
		4'd2: n_loc_oh_reg[161] = {13'd0, dist_reg[94], 2'd0};
		4'd3: n_loc_oh_reg[161] = {12'd0, dist_reg[94], 3'd0};
		4'd4: n_loc_oh_reg[161] = {11'd0, dist_reg[94], 4'd0};
		4'd5: n_loc_oh_reg[161] = {10'd0, dist_reg[94], 5'd0};
		4'd6: n_loc_oh_reg[161] = {9'd0, dist_reg[94], 6'd0};
		4'd7: n_loc_oh_reg[161] = {8'd0, dist_reg[94], 7'd0};
		4'd8: n_loc_oh_reg[161] = {7'd0, dist_reg[94], 8'd0};
		4'd9: n_loc_oh_reg[161] = {6'd0, dist_reg[94], 9'd0};
		4'd10: n_loc_oh_reg[161] = {5'd0, dist_reg[94], 10'd0};
		4'd11: n_loc_oh_reg[161] = {4'd0, dist_reg[94], 11'd0};
		4'd12: n_loc_oh_reg[161] = {3'd0, dist_reg[94], 12'd0};
		4'd13: n_loc_oh_reg[161] = {2'd0, dist_reg[94], 13'd0};
		4'd14: n_loc_oh_reg[161] = {1'd0, dist_reg[94], 14'd0};
		4'd15: n_loc_oh_reg[161] = {dist_reg[94], 15'd0};
	endcase
	case(loc_reg[162])
		4'd0: n_loc_oh_reg[162] = {15'd0, dist_reg[93]};
		4'd1: n_loc_oh_reg[162] = {14'd0, dist_reg[93], 1'd0};
		4'd2: n_loc_oh_reg[162] = {13'd0, dist_reg[93], 2'd0};
		4'd3: n_loc_oh_reg[162] = {12'd0, dist_reg[93], 3'd0};
		4'd4: n_loc_oh_reg[162] = {11'd0, dist_reg[93], 4'd0};
		4'd5: n_loc_oh_reg[162] = {10'd0, dist_reg[93], 5'd0};
		4'd6: n_loc_oh_reg[162] = {9'd0, dist_reg[93], 6'd0};
		4'd7: n_loc_oh_reg[162] = {8'd0, dist_reg[93], 7'd0};
		4'd8: n_loc_oh_reg[162] = {7'd0, dist_reg[93], 8'd0};
		4'd9: n_loc_oh_reg[162] = {6'd0, dist_reg[93], 9'd0};
		4'd10: n_loc_oh_reg[162] = {5'd0, dist_reg[93], 10'd0};
		4'd11: n_loc_oh_reg[162] = {4'd0, dist_reg[93], 11'd0};
		4'd12: n_loc_oh_reg[162] = {3'd0, dist_reg[93], 12'd0};
		4'd13: n_loc_oh_reg[162] = {2'd0, dist_reg[93], 13'd0};
		4'd14: n_loc_oh_reg[162] = {1'd0, dist_reg[93], 14'd0};
		4'd15: n_loc_oh_reg[162] = {dist_reg[93], 15'd0};
	endcase
	case(loc_reg[163])
		4'd0: n_loc_oh_reg[163] = {15'd0, dist_reg[92]};
		4'd1: n_loc_oh_reg[163] = {14'd0, dist_reg[92], 1'd0};
		4'd2: n_loc_oh_reg[163] = {13'd0, dist_reg[92], 2'd0};
		4'd3: n_loc_oh_reg[163] = {12'd0, dist_reg[92], 3'd0};
		4'd4: n_loc_oh_reg[163] = {11'd0, dist_reg[92], 4'd0};
		4'd5: n_loc_oh_reg[163] = {10'd0, dist_reg[92], 5'd0};
		4'd6: n_loc_oh_reg[163] = {9'd0, dist_reg[92], 6'd0};
		4'd7: n_loc_oh_reg[163] = {8'd0, dist_reg[92], 7'd0};
		4'd8: n_loc_oh_reg[163] = {7'd0, dist_reg[92], 8'd0};
		4'd9: n_loc_oh_reg[163] = {6'd0, dist_reg[92], 9'd0};
		4'd10: n_loc_oh_reg[163] = {5'd0, dist_reg[92], 10'd0};
		4'd11: n_loc_oh_reg[163] = {4'd0, dist_reg[92], 11'd0};
		4'd12: n_loc_oh_reg[163] = {3'd0, dist_reg[92], 12'd0};
		4'd13: n_loc_oh_reg[163] = {2'd0, dist_reg[92], 13'd0};
		4'd14: n_loc_oh_reg[163] = {1'd0, dist_reg[92], 14'd0};
		4'd15: n_loc_oh_reg[163] = {dist_reg[92], 15'd0};
	endcase
	case(loc_reg[164])
		4'd0: n_loc_oh_reg[164] = {15'd0, dist_reg[91]};
		4'd1: n_loc_oh_reg[164] = {14'd0, dist_reg[91], 1'd0};
		4'd2: n_loc_oh_reg[164] = {13'd0, dist_reg[91], 2'd0};
		4'd3: n_loc_oh_reg[164] = {12'd0, dist_reg[91], 3'd0};
		4'd4: n_loc_oh_reg[164] = {11'd0, dist_reg[91], 4'd0};
		4'd5: n_loc_oh_reg[164] = {10'd0, dist_reg[91], 5'd0};
		4'd6: n_loc_oh_reg[164] = {9'd0, dist_reg[91], 6'd0};
		4'd7: n_loc_oh_reg[164] = {8'd0, dist_reg[91], 7'd0};
		4'd8: n_loc_oh_reg[164] = {7'd0, dist_reg[91], 8'd0};
		4'd9: n_loc_oh_reg[164] = {6'd0, dist_reg[91], 9'd0};
		4'd10: n_loc_oh_reg[164] = {5'd0, dist_reg[91], 10'd0};
		4'd11: n_loc_oh_reg[164] = {4'd0, dist_reg[91], 11'd0};
		4'd12: n_loc_oh_reg[164] = {3'd0, dist_reg[91], 12'd0};
		4'd13: n_loc_oh_reg[164] = {2'd0, dist_reg[91], 13'd0};
		4'd14: n_loc_oh_reg[164] = {1'd0, dist_reg[91], 14'd0};
		4'd15: n_loc_oh_reg[164] = {dist_reg[91], 15'd0};
	endcase
	case(loc_reg[165])
		4'd0: n_loc_oh_reg[165] = {15'd0, dist_reg[90]};
		4'd1: n_loc_oh_reg[165] = {14'd0, dist_reg[90], 1'd0};
		4'd2: n_loc_oh_reg[165] = {13'd0, dist_reg[90], 2'd0};
		4'd3: n_loc_oh_reg[165] = {12'd0, dist_reg[90], 3'd0};
		4'd4: n_loc_oh_reg[165] = {11'd0, dist_reg[90], 4'd0};
		4'd5: n_loc_oh_reg[165] = {10'd0, dist_reg[90], 5'd0};
		4'd6: n_loc_oh_reg[165] = {9'd0, dist_reg[90], 6'd0};
		4'd7: n_loc_oh_reg[165] = {8'd0, dist_reg[90], 7'd0};
		4'd8: n_loc_oh_reg[165] = {7'd0, dist_reg[90], 8'd0};
		4'd9: n_loc_oh_reg[165] = {6'd0, dist_reg[90], 9'd0};
		4'd10: n_loc_oh_reg[165] = {5'd0, dist_reg[90], 10'd0};
		4'd11: n_loc_oh_reg[165] = {4'd0, dist_reg[90], 11'd0};
		4'd12: n_loc_oh_reg[165] = {3'd0, dist_reg[90], 12'd0};
		4'd13: n_loc_oh_reg[165] = {2'd0, dist_reg[90], 13'd0};
		4'd14: n_loc_oh_reg[165] = {1'd0, dist_reg[90], 14'd0};
		4'd15: n_loc_oh_reg[165] = {dist_reg[90], 15'd0};
	endcase
	case(loc_reg[166])
		4'd0: n_loc_oh_reg[166] = {15'd0, dist_reg[89]};
		4'd1: n_loc_oh_reg[166] = {14'd0, dist_reg[89], 1'd0};
		4'd2: n_loc_oh_reg[166] = {13'd0, dist_reg[89], 2'd0};
		4'd3: n_loc_oh_reg[166] = {12'd0, dist_reg[89], 3'd0};
		4'd4: n_loc_oh_reg[166] = {11'd0, dist_reg[89], 4'd0};
		4'd5: n_loc_oh_reg[166] = {10'd0, dist_reg[89], 5'd0};
		4'd6: n_loc_oh_reg[166] = {9'd0, dist_reg[89], 6'd0};
		4'd7: n_loc_oh_reg[166] = {8'd0, dist_reg[89], 7'd0};
		4'd8: n_loc_oh_reg[166] = {7'd0, dist_reg[89], 8'd0};
		4'd9: n_loc_oh_reg[166] = {6'd0, dist_reg[89], 9'd0};
		4'd10: n_loc_oh_reg[166] = {5'd0, dist_reg[89], 10'd0};
		4'd11: n_loc_oh_reg[166] = {4'd0, dist_reg[89], 11'd0};
		4'd12: n_loc_oh_reg[166] = {3'd0, dist_reg[89], 12'd0};
		4'd13: n_loc_oh_reg[166] = {2'd0, dist_reg[89], 13'd0};
		4'd14: n_loc_oh_reg[166] = {1'd0, dist_reg[89], 14'd0};
		4'd15: n_loc_oh_reg[166] = {dist_reg[89], 15'd0};
	endcase
	case(loc_reg[167])
		4'd0: n_loc_oh_reg[167] = {15'd0, dist_reg[88]};
		4'd1: n_loc_oh_reg[167] = {14'd0, dist_reg[88], 1'd0};
		4'd2: n_loc_oh_reg[167] = {13'd0, dist_reg[88], 2'd0};
		4'd3: n_loc_oh_reg[167] = {12'd0, dist_reg[88], 3'd0};
		4'd4: n_loc_oh_reg[167] = {11'd0, dist_reg[88], 4'd0};
		4'd5: n_loc_oh_reg[167] = {10'd0, dist_reg[88], 5'd0};
		4'd6: n_loc_oh_reg[167] = {9'd0, dist_reg[88], 6'd0};
		4'd7: n_loc_oh_reg[167] = {8'd0, dist_reg[88], 7'd0};
		4'd8: n_loc_oh_reg[167] = {7'd0, dist_reg[88], 8'd0};
		4'd9: n_loc_oh_reg[167] = {6'd0, dist_reg[88], 9'd0};
		4'd10: n_loc_oh_reg[167] = {5'd0, dist_reg[88], 10'd0};
		4'd11: n_loc_oh_reg[167] = {4'd0, dist_reg[88], 11'd0};
		4'd12: n_loc_oh_reg[167] = {3'd0, dist_reg[88], 12'd0};
		4'd13: n_loc_oh_reg[167] = {2'd0, dist_reg[88], 13'd0};
		4'd14: n_loc_oh_reg[167] = {1'd0, dist_reg[88], 14'd0};
		4'd15: n_loc_oh_reg[167] = {dist_reg[88], 15'd0};
	endcase
	case(loc_reg[168])
		4'd0: n_loc_oh_reg[168] = {15'd0, dist_reg[87]};
		4'd1: n_loc_oh_reg[168] = {14'd0, dist_reg[87], 1'd0};
		4'd2: n_loc_oh_reg[168] = {13'd0, dist_reg[87], 2'd0};
		4'd3: n_loc_oh_reg[168] = {12'd0, dist_reg[87], 3'd0};
		4'd4: n_loc_oh_reg[168] = {11'd0, dist_reg[87], 4'd0};
		4'd5: n_loc_oh_reg[168] = {10'd0, dist_reg[87], 5'd0};
		4'd6: n_loc_oh_reg[168] = {9'd0, dist_reg[87], 6'd0};
		4'd7: n_loc_oh_reg[168] = {8'd0, dist_reg[87], 7'd0};
		4'd8: n_loc_oh_reg[168] = {7'd0, dist_reg[87], 8'd0};
		4'd9: n_loc_oh_reg[168] = {6'd0, dist_reg[87], 9'd0};
		4'd10: n_loc_oh_reg[168] = {5'd0, dist_reg[87], 10'd0};
		4'd11: n_loc_oh_reg[168] = {4'd0, dist_reg[87], 11'd0};
		4'd12: n_loc_oh_reg[168] = {3'd0, dist_reg[87], 12'd0};
		4'd13: n_loc_oh_reg[168] = {2'd0, dist_reg[87], 13'd0};
		4'd14: n_loc_oh_reg[168] = {1'd0, dist_reg[87], 14'd0};
		4'd15: n_loc_oh_reg[168] = {dist_reg[87], 15'd0};
	endcase
	case(loc_reg[169])
		4'd0: n_loc_oh_reg[169] = {15'd0, dist_reg[86]};
		4'd1: n_loc_oh_reg[169] = {14'd0, dist_reg[86], 1'd0};
		4'd2: n_loc_oh_reg[169] = {13'd0, dist_reg[86], 2'd0};
		4'd3: n_loc_oh_reg[169] = {12'd0, dist_reg[86], 3'd0};
		4'd4: n_loc_oh_reg[169] = {11'd0, dist_reg[86], 4'd0};
		4'd5: n_loc_oh_reg[169] = {10'd0, dist_reg[86], 5'd0};
		4'd6: n_loc_oh_reg[169] = {9'd0, dist_reg[86], 6'd0};
		4'd7: n_loc_oh_reg[169] = {8'd0, dist_reg[86], 7'd0};
		4'd8: n_loc_oh_reg[169] = {7'd0, dist_reg[86], 8'd0};
		4'd9: n_loc_oh_reg[169] = {6'd0, dist_reg[86], 9'd0};
		4'd10: n_loc_oh_reg[169] = {5'd0, dist_reg[86], 10'd0};
		4'd11: n_loc_oh_reg[169] = {4'd0, dist_reg[86], 11'd0};
		4'd12: n_loc_oh_reg[169] = {3'd0, dist_reg[86], 12'd0};
		4'd13: n_loc_oh_reg[169] = {2'd0, dist_reg[86], 13'd0};
		4'd14: n_loc_oh_reg[169] = {1'd0, dist_reg[86], 14'd0};
		4'd15: n_loc_oh_reg[169] = {dist_reg[86], 15'd0};
	endcase
	case(loc_reg[170])
		4'd0: n_loc_oh_reg[170] = {15'd0, dist_reg[85]};
		4'd1: n_loc_oh_reg[170] = {14'd0, dist_reg[85], 1'd0};
		4'd2: n_loc_oh_reg[170] = {13'd0, dist_reg[85], 2'd0};
		4'd3: n_loc_oh_reg[170] = {12'd0, dist_reg[85], 3'd0};
		4'd4: n_loc_oh_reg[170] = {11'd0, dist_reg[85], 4'd0};
		4'd5: n_loc_oh_reg[170] = {10'd0, dist_reg[85], 5'd0};
		4'd6: n_loc_oh_reg[170] = {9'd0, dist_reg[85], 6'd0};
		4'd7: n_loc_oh_reg[170] = {8'd0, dist_reg[85], 7'd0};
		4'd8: n_loc_oh_reg[170] = {7'd0, dist_reg[85], 8'd0};
		4'd9: n_loc_oh_reg[170] = {6'd0, dist_reg[85], 9'd0};
		4'd10: n_loc_oh_reg[170] = {5'd0, dist_reg[85], 10'd0};
		4'd11: n_loc_oh_reg[170] = {4'd0, dist_reg[85], 11'd0};
		4'd12: n_loc_oh_reg[170] = {3'd0, dist_reg[85], 12'd0};
		4'd13: n_loc_oh_reg[170] = {2'd0, dist_reg[85], 13'd0};
		4'd14: n_loc_oh_reg[170] = {1'd0, dist_reg[85], 14'd0};
		4'd15: n_loc_oh_reg[170] = {dist_reg[85], 15'd0};
	endcase
	case(loc_reg[171])
		4'd0: n_loc_oh_reg[171] = {15'd0, dist_reg[84]};
		4'd1: n_loc_oh_reg[171] = {14'd0, dist_reg[84], 1'd0};
		4'd2: n_loc_oh_reg[171] = {13'd0, dist_reg[84], 2'd0};
		4'd3: n_loc_oh_reg[171] = {12'd0, dist_reg[84], 3'd0};
		4'd4: n_loc_oh_reg[171] = {11'd0, dist_reg[84], 4'd0};
		4'd5: n_loc_oh_reg[171] = {10'd0, dist_reg[84], 5'd0};
		4'd6: n_loc_oh_reg[171] = {9'd0, dist_reg[84], 6'd0};
		4'd7: n_loc_oh_reg[171] = {8'd0, dist_reg[84], 7'd0};
		4'd8: n_loc_oh_reg[171] = {7'd0, dist_reg[84], 8'd0};
		4'd9: n_loc_oh_reg[171] = {6'd0, dist_reg[84], 9'd0};
		4'd10: n_loc_oh_reg[171] = {5'd0, dist_reg[84], 10'd0};
		4'd11: n_loc_oh_reg[171] = {4'd0, dist_reg[84], 11'd0};
		4'd12: n_loc_oh_reg[171] = {3'd0, dist_reg[84], 12'd0};
		4'd13: n_loc_oh_reg[171] = {2'd0, dist_reg[84], 13'd0};
		4'd14: n_loc_oh_reg[171] = {1'd0, dist_reg[84], 14'd0};
		4'd15: n_loc_oh_reg[171] = {dist_reg[84], 15'd0};
	endcase
	case(loc_reg[172])
		4'd0: n_loc_oh_reg[172] = {15'd0, dist_reg[83]};
		4'd1: n_loc_oh_reg[172] = {14'd0, dist_reg[83], 1'd0};
		4'd2: n_loc_oh_reg[172] = {13'd0, dist_reg[83], 2'd0};
		4'd3: n_loc_oh_reg[172] = {12'd0, dist_reg[83], 3'd0};
		4'd4: n_loc_oh_reg[172] = {11'd0, dist_reg[83], 4'd0};
		4'd5: n_loc_oh_reg[172] = {10'd0, dist_reg[83], 5'd0};
		4'd6: n_loc_oh_reg[172] = {9'd0, dist_reg[83], 6'd0};
		4'd7: n_loc_oh_reg[172] = {8'd0, dist_reg[83], 7'd0};
		4'd8: n_loc_oh_reg[172] = {7'd0, dist_reg[83], 8'd0};
		4'd9: n_loc_oh_reg[172] = {6'd0, dist_reg[83], 9'd0};
		4'd10: n_loc_oh_reg[172] = {5'd0, dist_reg[83], 10'd0};
		4'd11: n_loc_oh_reg[172] = {4'd0, dist_reg[83], 11'd0};
		4'd12: n_loc_oh_reg[172] = {3'd0, dist_reg[83], 12'd0};
		4'd13: n_loc_oh_reg[172] = {2'd0, dist_reg[83], 13'd0};
		4'd14: n_loc_oh_reg[172] = {1'd0, dist_reg[83], 14'd0};
		4'd15: n_loc_oh_reg[172] = {dist_reg[83], 15'd0};
	endcase
	case(loc_reg[173])
		4'd0: n_loc_oh_reg[173] = {15'd0, dist_reg[82]};
		4'd1: n_loc_oh_reg[173] = {14'd0, dist_reg[82], 1'd0};
		4'd2: n_loc_oh_reg[173] = {13'd0, dist_reg[82], 2'd0};
		4'd3: n_loc_oh_reg[173] = {12'd0, dist_reg[82], 3'd0};
		4'd4: n_loc_oh_reg[173] = {11'd0, dist_reg[82], 4'd0};
		4'd5: n_loc_oh_reg[173] = {10'd0, dist_reg[82], 5'd0};
		4'd6: n_loc_oh_reg[173] = {9'd0, dist_reg[82], 6'd0};
		4'd7: n_loc_oh_reg[173] = {8'd0, dist_reg[82], 7'd0};
		4'd8: n_loc_oh_reg[173] = {7'd0, dist_reg[82], 8'd0};
		4'd9: n_loc_oh_reg[173] = {6'd0, dist_reg[82], 9'd0};
		4'd10: n_loc_oh_reg[173] = {5'd0, dist_reg[82], 10'd0};
		4'd11: n_loc_oh_reg[173] = {4'd0, dist_reg[82], 11'd0};
		4'd12: n_loc_oh_reg[173] = {3'd0, dist_reg[82], 12'd0};
		4'd13: n_loc_oh_reg[173] = {2'd0, dist_reg[82], 13'd0};
		4'd14: n_loc_oh_reg[173] = {1'd0, dist_reg[82], 14'd0};
		4'd15: n_loc_oh_reg[173] = {dist_reg[82], 15'd0};
	endcase
	case(loc_reg[174])
		4'd0: n_loc_oh_reg[174] = {15'd0, dist_reg[81]};
		4'd1: n_loc_oh_reg[174] = {14'd0, dist_reg[81], 1'd0};
		4'd2: n_loc_oh_reg[174] = {13'd0, dist_reg[81], 2'd0};
		4'd3: n_loc_oh_reg[174] = {12'd0, dist_reg[81], 3'd0};
		4'd4: n_loc_oh_reg[174] = {11'd0, dist_reg[81], 4'd0};
		4'd5: n_loc_oh_reg[174] = {10'd0, dist_reg[81], 5'd0};
		4'd6: n_loc_oh_reg[174] = {9'd0, dist_reg[81], 6'd0};
		4'd7: n_loc_oh_reg[174] = {8'd0, dist_reg[81], 7'd0};
		4'd8: n_loc_oh_reg[174] = {7'd0, dist_reg[81], 8'd0};
		4'd9: n_loc_oh_reg[174] = {6'd0, dist_reg[81], 9'd0};
		4'd10: n_loc_oh_reg[174] = {5'd0, dist_reg[81], 10'd0};
		4'd11: n_loc_oh_reg[174] = {4'd0, dist_reg[81], 11'd0};
		4'd12: n_loc_oh_reg[174] = {3'd0, dist_reg[81], 12'd0};
		4'd13: n_loc_oh_reg[174] = {2'd0, dist_reg[81], 13'd0};
		4'd14: n_loc_oh_reg[174] = {1'd0, dist_reg[81], 14'd0};
		4'd15: n_loc_oh_reg[174] = {dist_reg[81], 15'd0};
	endcase
	case(loc_reg[175])
		4'd0: n_loc_oh_reg[175] = {15'd0, dist_reg[80]};
		4'd1: n_loc_oh_reg[175] = {14'd0, dist_reg[80], 1'd0};
		4'd2: n_loc_oh_reg[175] = {13'd0, dist_reg[80], 2'd0};
		4'd3: n_loc_oh_reg[175] = {12'd0, dist_reg[80], 3'd0};
		4'd4: n_loc_oh_reg[175] = {11'd0, dist_reg[80], 4'd0};
		4'd5: n_loc_oh_reg[175] = {10'd0, dist_reg[80], 5'd0};
		4'd6: n_loc_oh_reg[175] = {9'd0, dist_reg[80], 6'd0};
		4'd7: n_loc_oh_reg[175] = {8'd0, dist_reg[80], 7'd0};
		4'd8: n_loc_oh_reg[175] = {7'd0, dist_reg[80], 8'd0};
		4'd9: n_loc_oh_reg[175] = {6'd0, dist_reg[80], 9'd0};
		4'd10: n_loc_oh_reg[175] = {5'd0, dist_reg[80], 10'd0};
		4'd11: n_loc_oh_reg[175] = {4'd0, dist_reg[80], 11'd0};
		4'd12: n_loc_oh_reg[175] = {3'd0, dist_reg[80], 12'd0};
		4'd13: n_loc_oh_reg[175] = {2'd0, dist_reg[80], 13'd0};
		4'd14: n_loc_oh_reg[175] = {1'd0, dist_reg[80], 14'd0};
		4'd15: n_loc_oh_reg[175] = {dist_reg[80], 15'd0};
	endcase
	case(loc_reg[176])
		4'd0: n_loc_oh_reg[176] = {15'd0, dist_reg[79]};
		4'd1: n_loc_oh_reg[176] = {14'd0, dist_reg[79], 1'd0};
		4'd2: n_loc_oh_reg[176] = {13'd0, dist_reg[79], 2'd0};
		4'd3: n_loc_oh_reg[176] = {12'd0, dist_reg[79], 3'd0};
		4'd4: n_loc_oh_reg[176] = {11'd0, dist_reg[79], 4'd0};
		4'd5: n_loc_oh_reg[176] = {10'd0, dist_reg[79], 5'd0};
		4'd6: n_loc_oh_reg[176] = {9'd0, dist_reg[79], 6'd0};
		4'd7: n_loc_oh_reg[176] = {8'd0, dist_reg[79], 7'd0};
		4'd8: n_loc_oh_reg[176] = {7'd0, dist_reg[79], 8'd0};
		4'd9: n_loc_oh_reg[176] = {6'd0, dist_reg[79], 9'd0};
		4'd10: n_loc_oh_reg[176] = {5'd0, dist_reg[79], 10'd0};
		4'd11: n_loc_oh_reg[176] = {4'd0, dist_reg[79], 11'd0};
		4'd12: n_loc_oh_reg[176] = {3'd0, dist_reg[79], 12'd0};
		4'd13: n_loc_oh_reg[176] = {2'd0, dist_reg[79], 13'd0};
		4'd14: n_loc_oh_reg[176] = {1'd0, dist_reg[79], 14'd0};
		4'd15: n_loc_oh_reg[176] = {dist_reg[79], 15'd0};
	endcase
	case(loc_reg[177])
		4'd0: n_loc_oh_reg[177] = {15'd0, dist_reg[78]};
		4'd1: n_loc_oh_reg[177] = {14'd0, dist_reg[78], 1'd0};
		4'd2: n_loc_oh_reg[177] = {13'd0, dist_reg[78], 2'd0};
		4'd3: n_loc_oh_reg[177] = {12'd0, dist_reg[78], 3'd0};
		4'd4: n_loc_oh_reg[177] = {11'd0, dist_reg[78], 4'd0};
		4'd5: n_loc_oh_reg[177] = {10'd0, dist_reg[78], 5'd0};
		4'd6: n_loc_oh_reg[177] = {9'd0, dist_reg[78], 6'd0};
		4'd7: n_loc_oh_reg[177] = {8'd0, dist_reg[78], 7'd0};
		4'd8: n_loc_oh_reg[177] = {7'd0, dist_reg[78], 8'd0};
		4'd9: n_loc_oh_reg[177] = {6'd0, dist_reg[78], 9'd0};
		4'd10: n_loc_oh_reg[177] = {5'd0, dist_reg[78], 10'd0};
		4'd11: n_loc_oh_reg[177] = {4'd0, dist_reg[78], 11'd0};
		4'd12: n_loc_oh_reg[177] = {3'd0, dist_reg[78], 12'd0};
		4'd13: n_loc_oh_reg[177] = {2'd0, dist_reg[78], 13'd0};
		4'd14: n_loc_oh_reg[177] = {1'd0, dist_reg[78], 14'd0};
		4'd15: n_loc_oh_reg[177] = {dist_reg[78], 15'd0};
	endcase
	case(loc_reg[178])
		4'd0: n_loc_oh_reg[178] = {15'd0, dist_reg[77]};
		4'd1: n_loc_oh_reg[178] = {14'd0, dist_reg[77], 1'd0};
		4'd2: n_loc_oh_reg[178] = {13'd0, dist_reg[77], 2'd0};
		4'd3: n_loc_oh_reg[178] = {12'd0, dist_reg[77], 3'd0};
		4'd4: n_loc_oh_reg[178] = {11'd0, dist_reg[77], 4'd0};
		4'd5: n_loc_oh_reg[178] = {10'd0, dist_reg[77], 5'd0};
		4'd6: n_loc_oh_reg[178] = {9'd0, dist_reg[77], 6'd0};
		4'd7: n_loc_oh_reg[178] = {8'd0, dist_reg[77], 7'd0};
		4'd8: n_loc_oh_reg[178] = {7'd0, dist_reg[77], 8'd0};
		4'd9: n_loc_oh_reg[178] = {6'd0, dist_reg[77], 9'd0};
		4'd10: n_loc_oh_reg[178] = {5'd0, dist_reg[77], 10'd0};
		4'd11: n_loc_oh_reg[178] = {4'd0, dist_reg[77], 11'd0};
		4'd12: n_loc_oh_reg[178] = {3'd0, dist_reg[77], 12'd0};
		4'd13: n_loc_oh_reg[178] = {2'd0, dist_reg[77], 13'd0};
		4'd14: n_loc_oh_reg[178] = {1'd0, dist_reg[77], 14'd0};
		4'd15: n_loc_oh_reg[178] = {dist_reg[77], 15'd0};
	endcase
	case(loc_reg[179])
		4'd0: n_loc_oh_reg[179] = {15'd0, dist_reg[76]};
		4'd1: n_loc_oh_reg[179] = {14'd0, dist_reg[76], 1'd0};
		4'd2: n_loc_oh_reg[179] = {13'd0, dist_reg[76], 2'd0};
		4'd3: n_loc_oh_reg[179] = {12'd0, dist_reg[76], 3'd0};
		4'd4: n_loc_oh_reg[179] = {11'd0, dist_reg[76], 4'd0};
		4'd5: n_loc_oh_reg[179] = {10'd0, dist_reg[76], 5'd0};
		4'd6: n_loc_oh_reg[179] = {9'd0, dist_reg[76], 6'd0};
		4'd7: n_loc_oh_reg[179] = {8'd0, dist_reg[76], 7'd0};
		4'd8: n_loc_oh_reg[179] = {7'd0, dist_reg[76], 8'd0};
		4'd9: n_loc_oh_reg[179] = {6'd0, dist_reg[76], 9'd0};
		4'd10: n_loc_oh_reg[179] = {5'd0, dist_reg[76], 10'd0};
		4'd11: n_loc_oh_reg[179] = {4'd0, dist_reg[76], 11'd0};
		4'd12: n_loc_oh_reg[179] = {3'd0, dist_reg[76], 12'd0};
		4'd13: n_loc_oh_reg[179] = {2'd0, dist_reg[76], 13'd0};
		4'd14: n_loc_oh_reg[179] = {1'd0, dist_reg[76], 14'd0};
		4'd15: n_loc_oh_reg[179] = {dist_reg[76], 15'd0};
	endcase
	case(loc_reg[180])
		4'd0: n_loc_oh_reg[180] = {15'd0, dist_reg[75]};
		4'd1: n_loc_oh_reg[180] = {14'd0, dist_reg[75], 1'd0};
		4'd2: n_loc_oh_reg[180] = {13'd0, dist_reg[75], 2'd0};
		4'd3: n_loc_oh_reg[180] = {12'd0, dist_reg[75], 3'd0};
		4'd4: n_loc_oh_reg[180] = {11'd0, dist_reg[75], 4'd0};
		4'd5: n_loc_oh_reg[180] = {10'd0, dist_reg[75], 5'd0};
		4'd6: n_loc_oh_reg[180] = {9'd0, dist_reg[75], 6'd0};
		4'd7: n_loc_oh_reg[180] = {8'd0, dist_reg[75], 7'd0};
		4'd8: n_loc_oh_reg[180] = {7'd0, dist_reg[75], 8'd0};
		4'd9: n_loc_oh_reg[180] = {6'd0, dist_reg[75], 9'd0};
		4'd10: n_loc_oh_reg[180] = {5'd0, dist_reg[75], 10'd0};
		4'd11: n_loc_oh_reg[180] = {4'd0, dist_reg[75], 11'd0};
		4'd12: n_loc_oh_reg[180] = {3'd0, dist_reg[75], 12'd0};
		4'd13: n_loc_oh_reg[180] = {2'd0, dist_reg[75], 13'd0};
		4'd14: n_loc_oh_reg[180] = {1'd0, dist_reg[75], 14'd0};
		4'd15: n_loc_oh_reg[180] = {dist_reg[75], 15'd0};
	endcase
	case(loc_reg[181])
		4'd0: n_loc_oh_reg[181] = {15'd0, dist_reg[74]};
		4'd1: n_loc_oh_reg[181] = {14'd0, dist_reg[74], 1'd0};
		4'd2: n_loc_oh_reg[181] = {13'd0, dist_reg[74], 2'd0};
		4'd3: n_loc_oh_reg[181] = {12'd0, dist_reg[74], 3'd0};
		4'd4: n_loc_oh_reg[181] = {11'd0, dist_reg[74], 4'd0};
		4'd5: n_loc_oh_reg[181] = {10'd0, dist_reg[74], 5'd0};
		4'd6: n_loc_oh_reg[181] = {9'd0, dist_reg[74], 6'd0};
		4'd7: n_loc_oh_reg[181] = {8'd0, dist_reg[74], 7'd0};
		4'd8: n_loc_oh_reg[181] = {7'd0, dist_reg[74], 8'd0};
		4'd9: n_loc_oh_reg[181] = {6'd0, dist_reg[74], 9'd0};
		4'd10: n_loc_oh_reg[181] = {5'd0, dist_reg[74], 10'd0};
		4'd11: n_loc_oh_reg[181] = {4'd0, dist_reg[74], 11'd0};
		4'd12: n_loc_oh_reg[181] = {3'd0, dist_reg[74], 12'd0};
		4'd13: n_loc_oh_reg[181] = {2'd0, dist_reg[74], 13'd0};
		4'd14: n_loc_oh_reg[181] = {1'd0, dist_reg[74], 14'd0};
		4'd15: n_loc_oh_reg[181] = {dist_reg[74], 15'd0};
	endcase
	case(loc_reg[182])
		4'd0: n_loc_oh_reg[182] = {15'd0, dist_reg[73]};
		4'd1: n_loc_oh_reg[182] = {14'd0, dist_reg[73], 1'd0};
		4'd2: n_loc_oh_reg[182] = {13'd0, dist_reg[73], 2'd0};
		4'd3: n_loc_oh_reg[182] = {12'd0, dist_reg[73], 3'd0};
		4'd4: n_loc_oh_reg[182] = {11'd0, dist_reg[73], 4'd0};
		4'd5: n_loc_oh_reg[182] = {10'd0, dist_reg[73], 5'd0};
		4'd6: n_loc_oh_reg[182] = {9'd0, dist_reg[73], 6'd0};
		4'd7: n_loc_oh_reg[182] = {8'd0, dist_reg[73], 7'd0};
		4'd8: n_loc_oh_reg[182] = {7'd0, dist_reg[73], 8'd0};
		4'd9: n_loc_oh_reg[182] = {6'd0, dist_reg[73], 9'd0};
		4'd10: n_loc_oh_reg[182] = {5'd0, dist_reg[73], 10'd0};
		4'd11: n_loc_oh_reg[182] = {4'd0, dist_reg[73], 11'd0};
		4'd12: n_loc_oh_reg[182] = {3'd0, dist_reg[73], 12'd0};
		4'd13: n_loc_oh_reg[182] = {2'd0, dist_reg[73], 13'd0};
		4'd14: n_loc_oh_reg[182] = {1'd0, dist_reg[73], 14'd0};
		4'd15: n_loc_oh_reg[182] = {dist_reg[73], 15'd0};
	endcase
	case(loc_reg[183])
		4'd0: n_loc_oh_reg[183] = {15'd0, dist_reg[72]};
		4'd1: n_loc_oh_reg[183] = {14'd0, dist_reg[72], 1'd0};
		4'd2: n_loc_oh_reg[183] = {13'd0, dist_reg[72], 2'd0};
		4'd3: n_loc_oh_reg[183] = {12'd0, dist_reg[72], 3'd0};
		4'd4: n_loc_oh_reg[183] = {11'd0, dist_reg[72], 4'd0};
		4'd5: n_loc_oh_reg[183] = {10'd0, dist_reg[72], 5'd0};
		4'd6: n_loc_oh_reg[183] = {9'd0, dist_reg[72], 6'd0};
		4'd7: n_loc_oh_reg[183] = {8'd0, dist_reg[72], 7'd0};
		4'd8: n_loc_oh_reg[183] = {7'd0, dist_reg[72], 8'd0};
		4'd9: n_loc_oh_reg[183] = {6'd0, dist_reg[72], 9'd0};
		4'd10: n_loc_oh_reg[183] = {5'd0, dist_reg[72], 10'd0};
		4'd11: n_loc_oh_reg[183] = {4'd0, dist_reg[72], 11'd0};
		4'd12: n_loc_oh_reg[183] = {3'd0, dist_reg[72], 12'd0};
		4'd13: n_loc_oh_reg[183] = {2'd0, dist_reg[72], 13'd0};
		4'd14: n_loc_oh_reg[183] = {1'd0, dist_reg[72], 14'd0};
		4'd15: n_loc_oh_reg[183] = {dist_reg[72], 15'd0};
	endcase
	case(loc_reg[184])
		4'd0: n_loc_oh_reg[184] = {15'd0, dist_reg[71]};
		4'd1: n_loc_oh_reg[184] = {14'd0, dist_reg[71], 1'd0};
		4'd2: n_loc_oh_reg[184] = {13'd0, dist_reg[71], 2'd0};
		4'd3: n_loc_oh_reg[184] = {12'd0, dist_reg[71], 3'd0};
		4'd4: n_loc_oh_reg[184] = {11'd0, dist_reg[71], 4'd0};
		4'd5: n_loc_oh_reg[184] = {10'd0, dist_reg[71], 5'd0};
		4'd6: n_loc_oh_reg[184] = {9'd0, dist_reg[71], 6'd0};
		4'd7: n_loc_oh_reg[184] = {8'd0, dist_reg[71], 7'd0};
		4'd8: n_loc_oh_reg[184] = {7'd0, dist_reg[71], 8'd0};
		4'd9: n_loc_oh_reg[184] = {6'd0, dist_reg[71], 9'd0};
		4'd10: n_loc_oh_reg[184] = {5'd0, dist_reg[71], 10'd0};
		4'd11: n_loc_oh_reg[184] = {4'd0, dist_reg[71], 11'd0};
		4'd12: n_loc_oh_reg[184] = {3'd0, dist_reg[71], 12'd0};
		4'd13: n_loc_oh_reg[184] = {2'd0, dist_reg[71], 13'd0};
		4'd14: n_loc_oh_reg[184] = {1'd0, dist_reg[71], 14'd0};
		4'd15: n_loc_oh_reg[184] = {dist_reg[71], 15'd0};
	endcase
	case(loc_reg[185])
		4'd0: n_loc_oh_reg[185] = {15'd0, dist_reg[70]};
		4'd1: n_loc_oh_reg[185] = {14'd0, dist_reg[70], 1'd0};
		4'd2: n_loc_oh_reg[185] = {13'd0, dist_reg[70], 2'd0};
		4'd3: n_loc_oh_reg[185] = {12'd0, dist_reg[70], 3'd0};
		4'd4: n_loc_oh_reg[185] = {11'd0, dist_reg[70], 4'd0};
		4'd5: n_loc_oh_reg[185] = {10'd0, dist_reg[70], 5'd0};
		4'd6: n_loc_oh_reg[185] = {9'd0, dist_reg[70], 6'd0};
		4'd7: n_loc_oh_reg[185] = {8'd0, dist_reg[70], 7'd0};
		4'd8: n_loc_oh_reg[185] = {7'd0, dist_reg[70], 8'd0};
		4'd9: n_loc_oh_reg[185] = {6'd0, dist_reg[70], 9'd0};
		4'd10: n_loc_oh_reg[185] = {5'd0, dist_reg[70], 10'd0};
		4'd11: n_loc_oh_reg[185] = {4'd0, dist_reg[70], 11'd0};
		4'd12: n_loc_oh_reg[185] = {3'd0, dist_reg[70], 12'd0};
		4'd13: n_loc_oh_reg[185] = {2'd0, dist_reg[70], 13'd0};
		4'd14: n_loc_oh_reg[185] = {1'd0, dist_reg[70], 14'd0};
		4'd15: n_loc_oh_reg[185] = {dist_reg[70], 15'd0};
	endcase
	case(loc_reg[186])
		4'd0: n_loc_oh_reg[186] = {15'd0, dist_reg[69]};
		4'd1: n_loc_oh_reg[186] = {14'd0, dist_reg[69], 1'd0};
		4'd2: n_loc_oh_reg[186] = {13'd0, dist_reg[69], 2'd0};
		4'd3: n_loc_oh_reg[186] = {12'd0, dist_reg[69], 3'd0};
		4'd4: n_loc_oh_reg[186] = {11'd0, dist_reg[69], 4'd0};
		4'd5: n_loc_oh_reg[186] = {10'd0, dist_reg[69], 5'd0};
		4'd6: n_loc_oh_reg[186] = {9'd0, dist_reg[69], 6'd0};
		4'd7: n_loc_oh_reg[186] = {8'd0, dist_reg[69], 7'd0};
		4'd8: n_loc_oh_reg[186] = {7'd0, dist_reg[69], 8'd0};
		4'd9: n_loc_oh_reg[186] = {6'd0, dist_reg[69], 9'd0};
		4'd10: n_loc_oh_reg[186] = {5'd0, dist_reg[69], 10'd0};
		4'd11: n_loc_oh_reg[186] = {4'd0, dist_reg[69], 11'd0};
		4'd12: n_loc_oh_reg[186] = {3'd0, dist_reg[69], 12'd0};
		4'd13: n_loc_oh_reg[186] = {2'd0, dist_reg[69], 13'd0};
		4'd14: n_loc_oh_reg[186] = {1'd0, dist_reg[69], 14'd0};
		4'd15: n_loc_oh_reg[186] = {dist_reg[69], 15'd0};
	endcase
	case(loc_reg[187])
		4'd0: n_loc_oh_reg[187] = {15'd0, dist_reg[68]};
		4'd1: n_loc_oh_reg[187] = {14'd0, dist_reg[68], 1'd0};
		4'd2: n_loc_oh_reg[187] = {13'd0, dist_reg[68], 2'd0};
		4'd3: n_loc_oh_reg[187] = {12'd0, dist_reg[68], 3'd0};
		4'd4: n_loc_oh_reg[187] = {11'd0, dist_reg[68], 4'd0};
		4'd5: n_loc_oh_reg[187] = {10'd0, dist_reg[68], 5'd0};
		4'd6: n_loc_oh_reg[187] = {9'd0, dist_reg[68], 6'd0};
		4'd7: n_loc_oh_reg[187] = {8'd0, dist_reg[68], 7'd0};
		4'd8: n_loc_oh_reg[187] = {7'd0, dist_reg[68], 8'd0};
		4'd9: n_loc_oh_reg[187] = {6'd0, dist_reg[68], 9'd0};
		4'd10: n_loc_oh_reg[187] = {5'd0, dist_reg[68], 10'd0};
		4'd11: n_loc_oh_reg[187] = {4'd0, dist_reg[68], 11'd0};
		4'd12: n_loc_oh_reg[187] = {3'd0, dist_reg[68], 12'd0};
		4'd13: n_loc_oh_reg[187] = {2'd0, dist_reg[68], 13'd0};
		4'd14: n_loc_oh_reg[187] = {1'd0, dist_reg[68], 14'd0};
		4'd15: n_loc_oh_reg[187] = {dist_reg[68], 15'd0};
	endcase
	case(loc_reg[188])
		4'd0: n_loc_oh_reg[188] = {15'd0, dist_reg[67]};
		4'd1: n_loc_oh_reg[188] = {14'd0, dist_reg[67], 1'd0};
		4'd2: n_loc_oh_reg[188] = {13'd0, dist_reg[67], 2'd0};
		4'd3: n_loc_oh_reg[188] = {12'd0, dist_reg[67], 3'd0};
		4'd4: n_loc_oh_reg[188] = {11'd0, dist_reg[67], 4'd0};
		4'd5: n_loc_oh_reg[188] = {10'd0, dist_reg[67], 5'd0};
		4'd6: n_loc_oh_reg[188] = {9'd0, dist_reg[67], 6'd0};
		4'd7: n_loc_oh_reg[188] = {8'd0, dist_reg[67], 7'd0};
		4'd8: n_loc_oh_reg[188] = {7'd0, dist_reg[67], 8'd0};
		4'd9: n_loc_oh_reg[188] = {6'd0, dist_reg[67], 9'd0};
		4'd10: n_loc_oh_reg[188] = {5'd0, dist_reg[67], 10'd0};
		4'd11: n_loc_oh_reg[188] = {4'd0, dist_reg[67], 11'd0};
		4'd12: n_loc_oh_reg[188] = {3'd0, dist_reg[67], 12'd0};
		4'd13: n_loc_oh_reg[188] = {2'd0, dist_reg[67], 13'd0};
		4'd14: n_loc_oh_reg[188] = {1'd0, dist_reg[67], 14'd0};
		4'd15: n_loc_oh_reg[188] = {dist_reg[67], 15'd0};
	endcase
	case(loc_reg[189])
		4'd0: n_loc_oh_reg[189] = {15'd0, dist_reg[66]};
		4'd1: n_loc_oh_reg[189] = {14'd0, dist_reg[66], 1'd0};
		4'd2: n_loc_oh_reg[189] = {13'd0, dist_reg[66], 2'd0};
		4'd3: n_loc_oh_reg[189] = {12'd0, dist_reg[66], 3'd0};
		4'd4: n_loc_oh_reg[189] = {11'd0, dist_reg[66], 4'd0};
		4'd5: n_loc_oh_reg[189] = {10'd0, dist_reg[66], 5'd0};
		4'd6: n_loc_oh_reg[189] = {9'd0, dist_reg[66], 6'd0};
		4'd7: n_loc_oh_reg[189] = {8'd0, dist_reg[66], 7'd0};
		4'd8: n_loc_oh_reg[189] = {7'd0, dist_reg[66], 8'd0};
		4'd9: n_loc_oh_reg[189] = {6'd0, dist_reg[66], 9'd0};
		4'd10: n_loc_oh_reg[189] = {5'd0, dist_reg[66], 10'd0};
		4'd11: n_loc_oh_reg[189] = {4'd0, dist_reg[66], 11'd0};
		4'd12: n_loc_oh_reg[189] = {3'd0, dist_reg[66], 12'd0};
		4'd13: n_loc_oh_reg[189] = {2'd0, dist_reg[66], 13'd0};
		4'd14: n_loc_oh_reg[189] = {1'd0, dist_reg[66], 14'd0};
		4'd15: n_loc_oh_reg[189] = {dist_reg[66], 15'd0};
	endcase
	case(loc_reg[190])
		4'd0: n_loc_oh_reg[190] = {15'd0, dist_reg[65]};
		4'd1: n_loc_oh_reg[190] = {14'd0, dist_reg[65], 1'd0};
		4'd2: n_loc_oh_reg[190] = {13'd0, dist_reg[65], 2'd0};
		4'd3: n_loc_oh_reg[190] = {12'd0, dist_reg[65], 3'd0};
		4'd4: n_loc_oh_reg[190] = {11'd0, dist_reg[65], 4'd0};
		4'd5: n_loc_oh_reg[190] = {10'd0, dist_reg[65], 5'd0};
		4'd6: n_loc_oh_reg[190] = {9'd0, dist_reg[65], 6'd0};
		4'd7: n_loc_oh_reg[190] = {8'd0, dist_reg[65], 7'd0};
		4'd8: n_loc_oh_reg[190] = {7'd0, dist_reg[65], 8'd0};
		4'd9: n_loc_oh_reg[190] = {6'd0, dist_reg[65], 9'd0};
		4'd10: n_loc_oh_reg[190] = {5'd0, dist_reg[65], 10'd0};
		4'd11: n_loc_oh_reg[190] = {4'd0, dist_reg[65], 11'd0};
		4'd12: n_loc_oh_reg[190] = {3'd0, dist_reg[65], 12'd0};
		4'd13: n_loc_oh_reg[190] = {2'd0, dist_reg[65], 13'd0};
		4'd14: n_loc_oh_reg[190] = {1'd0, dist_reg[65], 14'd0};
		4'd15: n_loc_oh_reg[190] = {dist_reg[65], 15'd0};
	endcase
	case(loc_reg[191])
		4'd0: n_loc_oh_reg[191] = {15'd0, dist_reg[64]};
		4'd1: n_loc_oh_reg[191] = {14'd0, dist_reg[64], 1'd0};
		4'd2: n_loc_oh_reg[191] = {13'd0, dist_reg[64], 2'd0};
		4'd3: n_loc_oh_reg[191] = {12'd0, dist_reg[64], 3'd0};
		4'd4: n_loc_oh_reg[191] = {11'd0, dist_reg[64], 4'd0};
		4'd5: n_loc_oh_reg[191] = {10'd0, dist_reg[64], 5'd0};
		4'd6: n_loc_oh_reg[191] = {9'd0, dist_reg[64], 6'd0};
		4'd7: n_loc_oh_reg[191] = {8'd0, dist_reg[64], 7'd0};
		4'd8: n_loc_oh_reg[191] = {7'd0, dist_reg[64], 8'd0};
		4'd9: n_loc_oh_reg[191] = {6'd0, dist_reg[64], 9'd0};
		4'd10: n_loc_oh_reg[191] = {5'd0, dist_reg[64], 10'd0};
		4'd11: n_loc_oh_reg[191] = {4'd0, dist_reg[64], 11'd0};
		4'd12: n_loc_oh_reg[191] = {3'd0, dist_reg[64], 12'd0};
		4'd13: n_loc_oh_reg[191] = {2'd0, dist_reg[64], 13'd0};
		4'd14: n_loc_oh_reg[191] = {1'd0, dist_reg[64], 14'd0};
		4'd15: n_loc_oh_reg[191] = {dist_reg[64], 15'd0};
	endcase
	case(loc_reg[192])
		4'd0: n_loc_oh_reg[192] = {15'd0, dist_reg[63]};
		4'd1: n_loc_oh_reg[192] = {14'd0, dist_reg[63], 1'd0};
		4'd2: n_loc_oh_reg[192] = {13'd0, dist_reg[63], 2'd0};
		4'd3: n_loc_oh_reg[192] = {12'd0, dist_reg[63], 3'd0};
		4'd4: n_loc_oh_reg[192] = {11'd0, dist_reg[63], 4'd0};
		4'd5: n_loc_oh_reg[192] = {10'd0, dist_reg[63], 5'd0};
		4'd6: n_loc_oh_reg[192] = {9'd0, dist_reg[63], 6'd0};
		4'd7: n_loc_oh_reg[192] = {8'd0, dist_reg[63], 7'd0};
		4'd8: n_loc_oh_reg[192] = {7'd0, dist_reg[63], 8'd0};
		4'd9: n_loc_oh_reg[192] = {6'd0, dist_reg[63], 9'd0};
		4'd10: n_loc_oh_reg[192] = {5'd0, dist_reg[63], 10'd0};
		4'd11: n_loc_oh_reg[192] = {4'd0, dist_reg[63], 11'd0};
		4'd12: n_loc_oh_reg[192] = {3'd0, dist_reg[63], 12'd0};
		4'd13: n_loc_oh_reg[192] = {2'd0, dist_reg[63], 13'd0};
		4'd14: n_loc_oh_reg[192] = {1'd0, dist_reg[63], 14'd0};
		4'd15: n_loc_oh_reg[192] = {dist_reg[63], 15'd0};
	endcase
	case(loc_reg[193])
		4'd0: n_loc_oh_reg[193] = {15'd0, dist_reg[62]};
		4'd1: n_loc_oh_reg[193] = {14'd0, dist_reg[62], 1'd0};
		4'd2: n_loc_oh_reg[193] = {13'd0, dist_reg[62], 2'd0};
		4'd3: n_loc_oh_reg[193] = {12'd0, dist_reg[62], 3'd0};
		4'd4: n_loc_oh_reg[193] = {11'd0, dist_reg[62], 4'd0};
		4'd5: n_loc_oh_reg[193] = {10'd0, dist_reg[62], 5'd0};
		4'd6: n_loc_oh_reg[193] = {9'd0, dist_reg[62], 6'd0};
		4'd7: n_loc_oh_reg[193] = {8'd0, dist_reg[62], 7'd0};
		4'd8: n_loc_oh_reg[193] = {7'd0, dist_reg[62], 8'd0};
		4'd9: n_loc_oh_reg[193] = {6'd0, dist_reg[62], 9'd0};
		4'd10: n_loc_oh_reg[193] = {5'd0, dist_reg[62], 10'd0};
		4'd11: n_loc_oh_reg[193] = {4'd0, dist_reg[62], 11'd0};
		4'd12: n_loc_oh_reg[193] = {3'd0, dist_reg[62], 12'd0};
		4'd13: n_loc_oh_reg[193] = {2'd0, dist_reg[62], 13'd0};
		4'd14: n_loc_oh_reg[193] = {1'd0, dist_reg[62], 14'd0};
		4'd15: n_loc_oh_reg[193] = {dist_reg[62], 15'd0};
	endcase
	case(loc_reg[194])
		4'd0: n_loc_oh_reg[194] = {15'd0, dist_reg[61]};
		4'd1: n_loc_oh_reg[194] = {14'd0, dist_reg[61], 1'd0};
		4'd2: n_loc_oh_reg[194] = {13'd0, dist_reg[61], 2'd0};
		4'd3: n_loc_oh_reg[194] = {12'd0, dist_reg[61], 3'd0};
		4'd4: n_loc_oh_reg[194] = {11'd0, dist_reg[61], 4'd0};
		4'd5: n_loc_oh_reg[194] = {10'd0, dist_reg[61], 5'd0};
		4'd6: n_loc_oh_reg[194] = {9'd0, dist_reg[61], 6'd0};
		4'd7: n_loc_oh_reg[194] = {8'd0, dist_reg[61], 7'd0};
		4'd8: n_loc_oh_reg[194] = {7'd0, dist_reg[61], 8'd0};
		4'd9: n_loc_oh_reg[194] = {6'd0, dist_reg[61], 9'd0};
		4'd10: n_loc_oh_reg[194] = {5'd0, dist_reg[61], 10'd0};
		4'd11: n_loc_oh_reg[194] = {4'd0, dist_reg[61], 11'd0};
		4'd12: n_loc_oh_reg[194] = {3'd0, dist_reg[61], 12'd0};
		4'd13: n_loc_oh_reg[194] = {2'd0, dist_reg[61], 13'd0};
		4'd14: n_loc_oh_reg[194] = {1'd0, dist_reg[61], 14'd0};
		4'd15: n_loc_oh_reg[194] = {dist_reg[61], 15'd0};
	endcase
	case(loc_reg[195])
		4'd0: n_loc_oh_reg[195] = {15'd0, dist_reg[60]};
		4'd1: n_loc_oh_reg[195] = {14'd0, dist_reg[60], 1'd0};
		4'd2: n_loc_oh_reg[195] = {13'd0, dist_reg[60], 2'd0};
		4'd3: n_loc_oh_reg[195] = {12'd0, dist_reg[60], 3'd0};
		4'd4: n_loc_oh_reg[195] = {11'd0, dist_reg[60], 4'd0};
		4'd5: n_loc_oh_reg[195] = {10'd0, dist_reg[60], 5'd0};
		4'd6: n_loc_oh_reg[195] = {9'd0, dist_reg[60], 6'd0};
		4'd7: n_loc_oh_reg[195] = {8'd0, dist_reg[60], 7'd0};
		4'd8: n_loc_oh_reg[195] = {7'd0, dist_reg[60], 8'd0};
		4'd9: n_loc_oh_reg[195] = {6'd0, dist_reg[60], 9'd0};
		4'd10: n_loc_oh_reg[195] = {5'd0, dist_reg[60], 10'd0};
		4'd11: n_loc_oh_reg[195] = {4'd0, dist_reg[60], 11'd0};
		4'd12: n_loc_oh_reg[195] = {3'd0, dist_reg[60], 12'd0};
		4'd13: n_loc_oh_reg[195] = {2'd0, dist_reg[60], 13'd0};
		4'd14: n_loc_oh_reg[195] = {1'd0, dist_reg[60], 14'd0};
		4'd15: n_loc_oh_reg[195] = {dist_reg[60], 15'd0};
	endcase
	case(loc_reg[196])
		4'd0: n_loc_oh_reg[196] = {15'd0, dist_reg[59]};
		4'd1: n_loc_oh_reg[196] = {14'd0, dist_reg[59], 1'd0};
		4'd2: n_loc_oh_reg[196] = {13'd0, dist_reg[59], 2'd0};
		4'd3: n_loc_oh_reg[196] = {12'd0, dist_reg[59], 3'd0};
		4'd4: n_loc_oh_reg[196] = {11'd0, dist_reg[59], 4'd0};
		4'd5: n_loc_oh_reg[196] = {10'd0, dist_reg[59], 5'd0};
		4'd6: n_loc_oh_reg[196] = {9'd0, dist_reg[59], 6'd0};
		4'd7: n_loc_oh_reg[196] = {8'd0, dist_reg[59], 7'd0};
		4'd8: n_loc_oh_reg[196] = {7'd0, dist_reg[59], 8'd0};
		4'd9: n_loc_oh_reg[196] = {6'd0, dist_reg[59], 9'd0};
		4'd10: n_loc_oh_reg[196] = {5'd0, dist_reg[59], 10'd0};
		4'd11: n_loc_oh_reg[196] = {4'd0, dist_reg[59], 11'd0};
		4'd12: n_loc_oh_reg[196] = {3'd0, dist_reg[59], 12'd0};
		4'd13: n_loc_oh_reg[196] = {2'd0, dist_reg[59], 13'd0};
		4'd14: n_loc_oh_reg[196] = {1'd0, dist_reg[59], 14'd0};
		4'd15: n_loc_oh_reg[196] = {dist_reg[59], 15'd0};
	endcase
	case(loc_reg[197])
		4'd0: n_loc_oh_reg[197] = {15'd0, dist_reg[58]};
		4'd1: n_loc_oh_reg[197] = {14'd0, dist_reg[58], 1'd0};
		4'd2: n_loc_oh_reg[197] = {13'd0, dist_reg[58], 2'd0};
		4'd3: n_loc_oh_reg[197] = {12'd0, dist_reg[58], 3'd0};
		4'd4: n_loc_oh_reg[197] = {11'd0, dist_reg[58], 4'd0};
		4'd5: n_loc_oh_reg[197] = {10'd0, dist_reg[58], 5'd0};
		4'd6: n_loc_oh_reg[197] = {9'd0, dist_reg[58], 6'd0};
		4'd7: n_loc_oh_reg[197] = {8'd0, dist_reg[58], 7'd0};
		4'd8: n_loc_oh_reg[197] = {7'd0, dist_reg[58], 8'd0};
		4'd9: n_loc_oh_reg[197] = {6'd0, dist_reg[58], 9'd0};
		4'd10: n_loc_oh_reg[197] = {5'd0, dist_reg[58], 10'd0};
		4'd11: n_loc_oh_reg[197] = {4'd0, dist_reg[58], 11'd0};
		4'd12: n_loc_oh_reg[197] = {3'd0, dist_reg[58], 12'd0};
		4'd13: n_loc_oh_reg[197] = {2'd0, dist_reg[58], 13'd0};
		4'd14: n_loc_oh_reg[197] = {1'd0, dist_reg[58], 14'd0};
		4'd15: n_loc_oh_reg[197] = {dist_reg[58], 15'd0};
	endcase
	case(loc_reg[198])
		4'd0: n_loc_oh_reg[198] = {15'd0, dist_reg[57]};
		4'd1: n_loc_oh_reg[198] = {14'd0, dist_reg[57], 1'd0};
		4'd2: n_loc_oh_reg[198] = {13'd0, dist_reg[57], 2'd0};
		4'd3: n_loc_oh_reg[198] = {12'd0, dist_reg[57], 3'd0};
		4'd4: n_loc_oh_reg[198] = {11'd0, dist_reg[57], 4'd0};
		4'd5: n_loc_oh_reg[198] = {10'd0, dist_reg[57], 5'd0};
		4'd6: n_loc_oh_reg[198] = {9'd0, dist_reg[57], 6'd0};
		4'd7: n_loc_oh_reg[198] = {8'd0, dist_reg[57], 7'd0};
		4'd8: n_loc_oh_reg[198] = {7'd0, dist_reg[57], 8'd0};
		4'd9: n_loc_oh_reg[198] = {6'd0, dist_reg[57], 9'd0};
		4'd10: n_loc_oh_reg[198] = {5'd0, dist_reg[57], 10'd0};
		4'd11: n_loc_oh_reg[198] = {4'd0, dist_reg[57], 11'd0};
		4'd12: n_loc_oh_reg[198] = {3'd0, dist_reg[57], 12'd0};
		4'd13: n_loc_oh_reg[198] = {2'd0, dist_reg[57], 13'd0};
		4'd14: n_loc_oh_reg[198] = {1'd0, dist_reg[57], 14'd0};
		4'd15: n_loc_oh_reg[198] = {dist_reg[57], 15'd0};
	endcase
	case(loc_reg[199])
		4'd0: n_loc_oh_reg[199] = {15'd0, dist_reg[56]};
		4'd1: n_loc_oh_reg[199] = {14'd0, dist_reg[56], 1'd0};
		4'd2: n_loc_oh_reg[199] = {13'd0, dist_reg[56], 2'd0};
		4'd3: n_loc_oh_reg[199] = {12'd0, dist_reg[56], 3'd0};
		4'd4: n_loc_oh_reg[199] = {11'd0, dist_reg[56], 4'd0};
		4'd5: n_loc_oh_reg[199] = {10'd0, dist_reg[56], 5'd0};
		4'd6: n_loc_oh_reg[199] = {9'd0, dist_reg[56], 6'd0};
		4'd7: n_loc_oh_reg[199] = {8'd0, dist_reg[56], 7'd0};
		4'd8: n_loc_oh_reg[199] = {7'd0, dist_reg[56], 8'd0};
		4'd9: n_loc_oh_reg[199] = {6'd0, dist_reg[56], 9'd0};
		4'd10: n_loc_oh_reg[199] = {5'd0, dist_reg[56], 10'd0};
		4'd11: n_loc_oh_reg[199] = {4'd0, dist_reg[56], 11'd0};
		4'd12: n_loc_oh_reg[199] = {3'd0, dist_reg[56], 12'd0};
		4'd13: n_loc_oh_reg[199] = {2'd0, dist_reg[56], 13'd0};
		4'd14: n_loc_oh_reg[199] = {1'd0, dist_reg[56], 14'd0};
		4'd15: n_loc_oh_reg[199] = {dist_reg[56], 15'd0};
	endcase
	case(loc_reg[200])
		4'd0: n_loc_oh_reg[200] = {15'd0, dist_reg[55]};
		4'd1: n_loc_oh_reg[200] = {14'd0, dist_reg[55], 1'd0};
		4'd2: n_loc_oh_reg[200] = {13'd0, dist_reg[55], 2'd0};
		4'd3: n_loc_oh_reg[200] = {12'd0, dist_reg[55], 3'd0};
		4'd4: n_loc_oh_reg[200] = {11'd0, dist_reg[55], 4'd0};
		4'd5: n_loc_oh_reg[200] = {10'd0, dist_reg[55], 5'd0};
		4'd6: n_loc_oh_reg[200] = {9'd0, dist_reg[55], 6'd0};
		4'd7: n_loc_oh_reg[200] = {8'd0, dist_reg[55], 7'd0};
		4'd8: n_loc_oh_reg[200] = {7'd0, dist_reg[55], 8'd0};
		4'd9: n_loc_oh_reg[200] = {6'd0, dist_reg[55], 9'd0};
		4'd10: n_loc_oh_reg[200] = {5'd0, dist_reg[55], 10'd0};
		4'd11: n_loc_oh_reg[200] = {4'd0, dist_reg[55], 11'd0};
		4'd12: n_loc_oh_reg[200] = {3'd0, dist_reg[55], 12'd0};
		4'd13: n_loc_oh_reg[200] = {2'd0, dist_reg[55], 13'd0};
		4'd14: n_loc_oh_reg[200] = {1'd0, dist_reg[55], 14'd0};
		4'd15: n_loc_oh_reg[200] = {dist_reg[55], 15'd0};
	endcase
	case(loc_reg[201])
		4'd0: n_loc_oh_reg[201] = {15'd0, dist_reg[54]};
		4'd1: n_loc_oh_reg[201] = {14'd0, dist_reg[54], 1'd0};
		4'd2: n_loc_oh_reg[201] = {13'd0, dist_reg[54], 2'd0};
		4'd3: n_loc_oh_reg[201] = {12'd0, dist_reg[54], 3'd0};
		4'd4: n_loc_oh_reg[201] = {11'd0, dist_reg[54], 4'd0};
		4'd5: n_loc_oh_reg[201] = {10'd0, dist_reg[54], 5'd0};
		4'd6: n_loc_oh_reg[201] = {9'd0, dist_reg[54], 6'd0};
		4'd7: n_loc_oh_reg[201] = {8'd0, dist_reg[54], 7'd0};
		4'd8: n_loc_oh_reg[201] = {7'd0, dist_reg[54], 8'd0};
		4'd9: n_loc_oh_reg[201] = {6'd0, dist_reg[54], 9'd0};
		4'd10: n_loc_oh_reg[201] = {5'd0, dist_reg[54], 10'd0};
		4'd11: n_loc_oh_reg[201] = {4'd0, dist_reg[54], 11'd0};
		4'd12: n_loc_oh_reg[201] = {3'd0, dist_reg[54], 12'd0};
		4'd13: n_loc_oh_reg[201] = {2'd0, dist_reg[54], 13'd0};
		4'd14: n_loc_oh_reg[201] = {1'd0, dist_reg[54], 14'd0};
		4'd15: n_loc_oh_reg[201] = {dist_reg[54], 15'd0};
	endcase
	case(loc_reg[202])
		4'd0: n_loc_oh_reg[202] = {15'd0, dist_reg[53]};
		4'd1: n_loc_oh_reg[202] = {14'd0, dist_reg[53], 1'd0};
		4'd2: n_loc_oh_reg[202] = {13'd0, dist_reg[53], 2'd0};
		4'd3: n_loc_oh_reg[202] = {12'd0, dist_reg[53], 3'd0};
		4'd4: n_loc_oh_reg[202] = {11'd0, dist_reg[53], 4'd0};
		4'd5: n_loc_oh_reg[202] = {10'd0, dist_reg[53], 5'd0};
		4'd6: n_loc_oh_reg[202] = {9'd0, dist_reg[53], 6'd0};
		4'd7: n_loc_oh_reg[202] = {8'd0, dist_reg[53], 7'd0};
		4'd8: n_loc_oh_reg[202] = {7'd0, dist_reg[53], 8'd0};
		4'd9: n_loc_oh_reg[202] = {6'd0, dist_reg[53], 9'd0};
		4'd10: n_loc_oh_reg[202] = {5'd0, dist_reg[53], 10'd0};
		4'd11: n_loc_oh_reg[202] = {4'd0, dist_reg[53], 11'd0};
		4'd12: n_loc_oh_reg[202] = {3'd0, dist_reg[53], 12'd0};
		4'd13: n_loc_oh_reg[202] = {2'd0, dist_reg[53], 13'd0};
		4'd14: n_loc_oh_reg[202] = {1'd0, dist_reg[53], 14'd0};
		4'd15: n_loc_oh_reg[202] = {dist_reg[53], 15'd0};
	endcase
	case(loc_reg[203])
		4'd0: n_loc_oh_reg[203] = {15'd0, dist_reg[52]};
		4'd1: n_loc_oh_reg[203] = {14'd0, dist_reg[52], 1'd0};
		4'd2: n_loc_oh_reg[203] = {13'd0, dist_reg[52], 2'd0};
		4'd3: n_loc_oh_reg[203] = {12'd0, dist_reg[52], 3'd0};
		4'd4: n_loc_oh_reg[203] = {11'd0, dist_reg[52], 4'd0};
		4'd5: n_loc_oh_reg[203] = {10'd0, dist_reg[52], 5'd0};
		4'd6: n_loc_oh_reg[203] = {9'd0, dist_reg[52], 6'd0};
		4'd7: n_loc_oh_reg[203] = {8'd0, dist_reg[52], 7'd0};
		4'd8: n_loc_oh_reg[203] = {7'd0, dist_reg[52], 8'd0};
		4'd9: n_loc_oh_reg[203] = {6'd0, dist_reg[52], 9'd0};
		4'd10: n_loc_oh_reg[203] = {5'd0, dist_reg[52], 10'd0};
		4'd11: n_loc_oh_reg[203] = {4'd0, dist_reg[52], 11'd0};
		4'd12: n_loc_oh_reg[203] = {3'd0, dist_reg[52], 12'd0};
		4'd13: n_loc_oh_reg[203] = {2'd0, dist_reg[52], 13'd0};
		4'd14: n_loc_oh_reg[203] = {1'd0, dist_reg[52], 14'd0};
		4'd15: n_loc_oh_reg[203] = {dist_reg[52], 15'd0};
	endcase
	case(loc_reg[204])
		4'd0: n_loc_oh_reg[204] = {15'd0, dist_reg[51]};
		4'd1: n_loc_oh_reg[204] = {14'd0, dist_reg[51], 1'd0};
		4'd2: n_loc_oh_reg[204] = {13'd0, dist_reg[51], 2'd0};
		4'd3: n_loc_oh_reg[204] = {12'd0, dist_reg[51], 3'd0};
		4'd4: n_loc_oh_reg[204] = {11'd0, dist_reg[51], 4'd0};
		4'd5: n_loc_oh_reg[204] = {10'd0, dist_reg[51], 5'd0};
		4'd6: n_loc_oh_reg[204] = {9'd0, dist_reg[51], 6'd0};
		4'd7: n_loc_oh_reg[204] = {8'd0, dist_reg[51], 7'd0};
		4'd8: n_loc_oh_reg[204] = {7'd0, dist_reg[51], 8'd0};
		4'd9: n_loc_oh_reg[204] = {6'd0, dist_reg[51], 9'd0};
		4'd10: n_loc_oh_reg[204] = {5'd0, dist_reg[51], 10'd0};
		4'd11: n_loc_oh_reg[204] = {4'd0, dist_reg[51], 11'd0};
		4'd12: n_loc_oh_reg[204] = {3'd0, dist_reg[51], 12'd0};
		4'd13: n_loc_oh_reg[204] = {2'd0, dist_reg[51], 13'd0};
		4'd14: n_loc_oh_reg[204] = {1'd0, dist_reg[51], 14'd0};
		4'd15: n_loc_oh_reg[204] = {dist_reg[51], 15'd0};
	endcase
	case(loc_reg[205])
		4'd0: n_loc_oh_reg[205] = {15'd0, dist_reg[50]};
		4'd1: n_loc_oh_reg[205] = {14'd0, dist_reg[50], 1'd0};
		4'd2: n_loc_oh_reg[205] = {13'd0, dist_reg[50], 2'd0};
		4'd3: n_loc_oh_reg[205] = {12'd0, dist_reg[50], 3'd0};
		4'd4: n_loc_oh_reg[205] = {11'd0, dist_reg[50], 4'd0};
		4'd5: n_loc_oh_reg[205] = {10'd0, dist_reg[50], 5'd0};
		4'd6: n_loc_oh_reg[205] = {9'd0, dist_reg[50], 6'd0};
		4'd7: n_loc_oh_reg[205] = {8'd0, dist_reg[50], 7'd0};
		4'd8: n_loc_oh_reg[205] = {7'd0, dist_reg[50], 8'd0};
		4'd9: n_loc_oh_reg[205] = {6'd0, dist_reg[50], 9'd0};
		4'd10: n_loc_oh_reg[205] = {5'd0, dist_reg[50], 10'd0};
		4'd11: n_loc_oh_reg[205] = {4'd0, dist_reg[50], 11'd0};
		4'd12: n_loc_oh_reg[205] = {3'd0, dist_reg[50], 12'd0};
		4'd13: n_loc_oh_reg[205] = {2'd0, dist_reg[50], 13'd0};
		4'd14: n_loc_oh_reg[205] = {1'd0, dist_reg[50], 14'd0};
		4'd15: n_loc_oh_reg[205] = {dist_reg[50], 15'd0};
	endcase
	case(loc_reg[206])
		4'd0: n_loc_oh_reg[206] = {15'd0, dist_reg[49]};
		4'd1: n_loc_oh_reg[206] = {14'd0, dist_reg[49], 1'd0};
		4'd2: n_loc_oh_reg[206] = {13'd0, dist_reg[49], 2'd0};
		4'd3: n_loc_oh_reg[206] = {12'd0, dist_reg[49], 3'd0};
		4'd4: n_loc_oh_reg[206] = {11'd0, dist_reg[49], 4'd0};
		4'd5: n_loc_oh_reg[206] = {10'd0, dist_reg[49], 5'd0};
		4'd6: n_loc_oh_reg[206] = {9'd0, dist_reg[49], 6'd0};
		4'd7: n_loc_oh_reg[206] = {8'd0, dist_reg[49], 7'd0};
		4'd8: n_loc_oh_reg[206] = {7'd0, dist_reg[49], 8'd0};
		4'd9: n_loc_oh_reg[206] = {6'd0, dist_reg[49], 9'd0};
		4'd10: n_loc_oh_reg[206] = {5'd0, dist_reg[49], 10'd0};
		4'd11: n_loc_oh_reg[206] = {4'd0, dist_reg[49], 11'd0};
		4'd12: n_loc_oh_reg[206] = {3'd0, dist_reg[49], 12'd0};
		4'd13: n_loc_oh_reg[206] = {2'd0, dist_reg[49], 13'd0};
		4'd14: n_loc_oh_reg[206] = {1'd0, dist_reg[49], 14'd0};
		4'd15: n_loc_oh_reg[206] = {dist_reg[49], 15'd0};
	endcase
	case(loc_reg[207])
		4'd0: n_loc_oh_reg[207] = {15'd0, dist_reg[48]};
		4'd1: n_loc_oh_reg[207] = {14'd0, dist_reg[48], 1'd0};
		4'd2: n_loc_oh_reg[207] = {13'd0, dist_reg[48], 2'd0};
		4'd3: n_loc_oh_reg[207] = {12'd0, dist_reg[48], 3'd0};
		4'd4: n_loc_oh_reg[207] = {11'd0, dist_reg[48], 4'd0};
		4'd5: n_loc_oh_reg[207] = {10'd0, dist_reg[48], 5'd0};
		4'd6: n_loc_oh_reg[207] = {9'd0, dist_reg[48], 6'd0};
		4'd7: n_loc_oh_reg[207] = {8'd0, dist_reg[48], 7'd0};
		4'd8: n_loc_oh_reg[207] = {7'd0, dist_reg[48], 8'd0};
		4'd9: n_loc_oh_reg[207] = {6'd0, dist_reg[48], 9'd0};
		4'd10: n_loc_oh_reg[207] = {5'd0, dist_reg[48], 10'd0};
		4'd11: n_loc_oh_reg[207] = {4'd0, dist_reg[48], 11'd0};
		4'd12: n_loc_oh_reg[207] = {3'd0, dist_reg[48], 12'd0};
		4'd13: n_loc_oh_reg[207] = {2'd0, dist_reg[48], 13'd0};
		4'd14: n_loc_oh_reg[207] = {1'd0, dist_reg[48], 14'd0};
		4'd15: n_loc_oh_reg[207] = {dist_reg[48], 15'd0};
	endcase
	case(loc_reg[208])
		4'd0: n_loc_oh_reg[208] = {15'd0, dist_reg[47]};
		4'd1: n_loc_oh_reg[208] = {14'd0, dist_reg[47], 1'd0};
		4'd2: n_loc_oh_reg[208] = {13'd0, dist_reg[47], 2'd0};
		4'd3: n_loc_oh_reg[208] = {12'd0, dist_reg[47], 3'd0};
		4'd4: n_loc_oh_reg[208] = {11'd0, dist_reg[47], 4'd0};
		4'd5: n_loc_oh_reg[208] = {10'd0, dist_reg[47], 5'd0};
		4'd6: n_loc_oh_reg[208] = {9'd0, dist_reg[47], 6'd0};
		4'd7: n_loc_oh_reg[208] = {8'd0, dist_reg[47], 7'd0};
		4'd8: n_loc_oh_reg[208] = {7'd0, dist_reg[47], 8'd0};
		4'd9: n_loc_oh_reg[208] = {6'd0, dist_reg[47], 9'd0};
		4'd10: n_loc_oh_reg[208] = {5'd0, dist_reg[47], 10'd0};
		4'd11: n_loc_oh_reg[208] = {4'd0, dist_reg[47], 11'd0};
		4'd12: n_loc_oh_reg[208] = {3'd0, dist_reg[47], 12'd0};
		4'd13: n_loc_oh_reg[208] = {2'd0, dist_reg[47], 13'd0};
		4'd14: n_loc_oh_reg[208] = {1'd0, dist_reg[47], 14'd0};
		4'd15: n_loc_oh_reg[208] = {dist_reg[47], 15'd0};
	endcase
	case(loc_reg[209])
		4'd0: n_loc_oh_reg[209] = {15'd0, dist_reg[46]};
		4'd1: n_loc_oh_reg[209] = {14'd0, dist_reg[46], 1'd0};
		4'd2: n_loc_oh_reg[209] = {13'd0, dist_reg[46], 2'd0};
		4'd3: n_loc_oh_reg[209] = {12'd0, dist_reg[46], 3'd0};
		4'd4: n_loc_oh_reg[209] = {11'd0, dist_reg[46], 4'd0};
		4'd5: n_loc_oh_reg[209] = {10'd0, dist_reg[46], 5'd0};
		4'd6: n_loc_oh_reg[209] = {9'd0, dist_reg[46], 6'd0};
		4'd7: n_loc_oh_reg[209] = {8'd0, dist_reg[46], 7'd0};
		4'd8: n_loc_oh_reg[209] = {7'd0, dist_reg[46], 8'd0};
		4'd9: n_loc_oh_reg[209] = {6'd0, dist_reg[46], 9'd0};
		4'd10: n_loc_oh_reg[209] = {5'd0, dist_reg[46], 10'd0};
		4'd11: n_loc_oh_reg[209] = {4'd0, dist_reg[46], 11'd0};
		4'd12: n_loc_oh_reg[209] = {3'd0, dist_reg[46], 12'd0};
		4'd13: n_loc_oh_reg[209] = {2'd0, dist_reg[46], 13'd0};
		4'd14: n_loc_oh_reg[209] = {1'd0, dist_reg[46], 14'd0};
		4'd15: n_loc_oh_reg[209] = {dist_reg[46], 15'd0};
	endcase
	case(loc_reg[210])
		4'd0: n_loc_oh_reg[210] = {15'd0, dist_reg[45]};
		4'd1: n_loc_oh_reg[210] = {14'd0, dist_reg[45], 1'd0};
		4'd2: n_loc_oh_reg[210] = {13'd0, dist_reg[45], 2'd0};
		4'd3: n_loc_oh_reg[210] = {12'd0, dist_reg[45], 3'd0};
		4'd4: n_loc_oh_reg[210] = {11'd0, dist_reg[45], 4'd0};
		4'd5: n_loc_oh_reg[210] = {10'd0, dist_reg[45], 5'd0};
		4'd6: n_loc_oh_reg[210] = {9'd0, dist_reg[45], 6'd0};
		4'd7: n_loc_oh_reg[210] = {8'd0, dist_reg[45], 7'd0};
		4'd8: n_loc_oh_reg[210] = {7'd0, dist_reg[45], 8'd0};
		4'd9: n_loc_oh_reg[210] = {6'd0, dist_reg[45], 9'd0};
		4'd10: n_loc_oh_reg[210] = {5'd0, dist_reg[45], 10'd0};
		4'd11: n_loc_oh_reg[210] = {4'd0, dist_reg[45], 11'd0};
		4'd12: n_loc_oh_reg[210] = {3'd0, dist_reg[45], 12'd0};
		4'd13: n_loc_oh_reg[210] = {2'd0, dist_reg[45], 13'd0};
		4'd14: n_loc_oh_reg[210] = {1'd0, dist_reg[45], 14'd0};
		4'd15: n_loc_oh_reg[210] = {dist_reg[45], 15'd0};
	endcase
	case(loc_reg[211])
		4'd0: n_loc_oh_reg[211] = {15'd0, dist_reg[44]};
		4'd1: n_loc_oh_reg[211] = {14'd0, dist_reg[44], 1'd0};
		4'd2: n_loc_oh_reg[211] = {13'd0, dist_reg[44], 2'd0};
		4'd3: n_loc_oh_reg[211] = {12'd0, dist_reg[44], 3'd0};
		4'd4: n_loc_oh_reg[211] = {11'd0, dist_reg[44], 4'd0};
		4'd5: n_loc_oh_reg[211] = {10'd0, dist_reg[44], 5'd0};
		4'd6: n_loc_oh_reg[211] = {9'd0, dist_reg[44], 6'd0};
		4'd7: n_loc_oh_reg[211] = {8'd0, dist_reg[44], 7'd0};
		4'd8: n_loc_oh_reg[211] = {7'd0, dist_reg[44], 8'd0};
		4'd9: n_loc_oh_reg[211] = {6'd0, dist_reg[44], 9'd0};
		4'd10: n_loc_oh_reg[211] = {5'd0, dist_reg[44], 10'd0};
		4'd11: n_loc_oh_reg[211] = {4'd0, dist_reg[44], 11'd0};
		4'd12: n_loc_oh_reg[211] = {3'd0, dist_reg[44], 12'd0};
		4'd13: n_loc_oh_reg[211] = {2'd0, dist_reg[44], 13'd0};
		4'd14: n_loc_oh_reg[211] = {1'd0, dist_reg[44], 14'd0};
		4'd15: n_loc_oh_reg[211] = {dist_reg[44], 15'd0};
	endcase
	case(loc_reg[212])
		4'd0: n_loc_oh_reg[212] = {15'd0, dist_reg[43]};
		4'd1: n_loc_oh_reg[212] = {14'd0, dist_reg[43], 1'd0};
		4'd2: n_loc_oh_reg[212] = {13'd0, dist_reg[43], 2'd0};
		4'd3: n_loc_oh_reg[212] = {12'd0, dist_reg[43], 3'd0};
		4'd4: n_loc_oh_reg[212] = {11'd0, dist_reg[43], 4'd0};
		4'd5: n_loc_oh_reg[212] = {10'd0, dist_reg[43], 5'd0};
		4'd6: n_loc_oh_reg[212] = {9'd0, dist_reg[43], 6'd0};
		4'd7: n_loc_oh_reg[212] = {8'd0, dist_reg[43], 7'd0};
		4'd8: n_loc_oh_reg[212] = {7'd0, dist_reg[43], 8'd0};
		4'd9: n_loc_oh_reg[212] = {6'd0, dist_reg[43], 9'd0};
		4'd10: n_loc_oh_reg[212] = {5'd0, dist_reg[43], 10'd0};
		4'd11: n_loc_oh_reg[212] = {4'd0, dist_reg[43], 11'd0};
		4'd12: n_loc_oh_reg[212] = {3'd0, dist_reg[43], 12'd0};
		4'd13: n_loc_oh_reg[212] = {2'd0, dist_reg[43], 13'd0};
		4'd14: n_loc_oh_reg[212] = {1'd0, dist_reg[43], 14'd0};
		4'd15: n_loc_oh_reg[212] = {dist_reg[43], 15'd0};
	endcase
	case(loc_reg[213])
		4'd0: n_loc_oh_reg[213] = {15'd0, dist_reg[42]};
		4'd1: n_loc_oh_reg[213] = {14'd0, dist_reg[42], 1'd0};
		4'd2: n_loc_oh_reg[213] = {13'd0, dist_reg[42], 2'd0};
		4'd3: n_loc_oh_reg[213] = {12'd0, dist_reg[42], 3'd0};
		4'd4: n_loc_oh_reg[213] = {11'd0, dist_reg[42], 4'd0};
		4'd5: n_loc_oh_reg[213] = {10'd0, dist_reg[42], 5'd0};
		4'd6: n_loc_oh_reg[213] = {9'd0, dist_reg[42], 6'd0};
		4'd7: n_loc_oh_reg[213] = {8'd0, dist_reg[42], 7'd0};
		4'd8: n_loc_oh_reg[213] = {7'd0, dist_reg[42], 8'd0};
		4'd9: n_loc_oh_reg[213] = {6'd0, dist_reg[42], 9'd0};
		4'd10: n_loc_oh_reg[213] = {5'd0, dist_reg[42], 10'd0};
		4'd11: n_loc_oh_reg[213] = {4'd0, dist_reg[42], 11'd0};
		4'd12: n_loc_oh_reg[213] = {3'd0, dist_reg[42], 12'd0};
		4'd13: n_loc_oh_reg[213] = {2'd0, dist_reg[42], 13'd0};
		4'd14: n_loc_oh_reg[213] = {1'd0, dist_reg[42], 14'd0};
		4'd15: n_loc_oh_reg[213] = {dist_reg[42], 15'd0};
	endcase
	case(loc_reg[214])
		4'd0: n_loc_oh_reg[214] = {15'd0, dist_reg[41]};
		4'd1: n_loc_oh_reg[214] = {14'd0, dist_reg[41], 1'd0};
		4'd2: n_loc_oh_reg[214] = {13'd0, dist_reg[41], 2'd0};
		4'd3: n_loc_oh_reg[214] = {12'd0, dist_reg[41], 3'd0};
		4'd4: n_loc_oh_reg[214] = {11'd0, dist_reg[41], 4'd0};
		4'd5: n_loc_oh_reg[214] = {10'd0, dist_reg[41], 5'd0};
		4'd6: n_loc_oh_reg[214] = {9'd0, dist_reg[41], 6'd0};
		4'd7: n_loc_oh_reg[214] = {8'd0, dist_reg[41], 7'd0};
		4'd8: n_loc_oh_reg[214] = {7'd0, dist_reg[41], 8'd0};
		4'd9: n_loc_oh_reg[214] = {6'd0, dist_reg[41], 9'd0};
		4'd10: n_loc_oh_reg[214] = {5'd0, dist_reg[41], 10'd0};
		4'd11: n_loc_oh_reg[214] = {4'd0, dist_reg[41], 11'd0};
		4'd12: n_loc_oh_reg[214] = {3'd0, dist_reg[41], 12'd0};
		4'd13: n_loc_oh_reg[214] = {2'd0, dist_reg[41], 13'd0};
		4'd14: n_loc_oh_reg[214] = {1'd0, dist_reg[41], 14'd0};
		4'd15: n_loc_oh_reg[214] = {dist_reg[41], 15'd0};
	endcase
	case(loc_reg[215])
		4'd0: n_loc_oh_reg[215] = {15'd0, dist_reg[40]};
		4'd1: n_loc_oh_reg[215] = {14'd0, dist_reg[40], 1'd0};
		4'd2: n_loc_oh_reg[215] = {13'd0, dist_reg[40], 2'd0};
		4'd3: n_loc_oh_reg[215] = {12'd0, dist_reg[40], 3'd0};
		4'd4: n_loc_oh_reg[215] = {11'd0, dist_reg[40], 4'd0};
		4'd5: n_loc_oh_reg[215] = {10'd0, dist_reg[40], 5'd0};
		4'd6: n_loc_oh_reg[215] = {9'd0, dist_reg[40], 6'd0};
		4'd7: n_loc_oh_reg[215] = {8'd0, dist_reg[40], 7'd0};
		4'd8: n_loc_oh_reg[215] = {7'd0, dist_reg[40], 8'd0};
		4'd9: n_loc_oh_reg[215] = {6'd0, dist_reg[40], 9'd0};
		4'd10: n_loc_oh_reg[215] = {5'd0, dist_reg[40], 10'd0};
		4'd11: n_loc_oh_reg[215] = {4'd0, dist_reg[40], 11'd0};
		4'd12: n_loc_oh_reg[215] = {3'd0, dist_reg[40], 12'd0};
		4'd13: n_loc_oh_reg[215] = {2'd0, dist_reg[40], 13'd0};
		4'd14: n_loc_oh_reg[215] = {1'd0, dist_reg[40], 14'd0};
		4'd15: n_loc_oh_reg[215] = {dist_reg[40], 15'd0};
	endcase
	case(loc_reg[216])
		4'd0: n_loc_oh_reg[216] = {15'd0, dist_reg[39]};
		4'd1: n_loc_oh_reg[216] = {14'd0, dist_reg[39], 1'd0};
		4'd2: n_loc_oh_reg[216] = {13'd0, dist_reg[39], 2'd0};
		4'd3: n_loc_oh_reg[216] = {12'd0, dist_reg[39], 3'd0};
		4'd4: n_loc_oh_reg[216] = {11'd0, dist_reg[39], 4'd0};
		4'd5: n_loc_oh_reg[216] = {10'd0, dist_reg[39], 5'd0};
		4'd6: n_loc_oh_reg[216] = {9'd0, dist_reg[39], 6'd0};
		4'd7: n_loc_oh_reg[216] = {8'd0, dist_reg[39], 7'd0};
		4'd8: n_loc_oh_reg[216] = {7'd0, dist_reg[39], 8'd0};
		4'd9: n_loc_oh_reg[216] = {6'd0, dist_reg[39], 9'd0};
		4'd10: n_loc_oh_reg[216] = {5'd0, dist_reg[39], 10'd0};
		4'd11: n_loc_oh_reg[216] = {4'd0, dist_reg[39], 11'd0};
		4'd12: n_loc_oh_reg[216] = {3'd0, dist_reg[39], 12'd0};
		4'd13: n_loc_oh_reg[216] = {2'd0, dist_reg[39], 13'd0};
		4'd14: n_loc_oh_reg[216] = {1'd0, dist_reg[39], 14'd0};
		4'd15: n_loc_oh_reg[216] = {dist_reg[39], 15'd0};
	endcase
	case(loc_reg[217])
		4'd0: n_loc_oh_reg[217] = {15'd0, dist_reg[38]};
		4'd1: n_loc_oh_reg[217] = {14'd0, dist_reg[38], 1'd0};
		4'd2: n_loc_oh_reg[217] = {13'd0, dist_reg[38], 2'd0};
		4'd3: n_loc_oh_reg[217] = {12'd0, dist_reg[38], 3'd0};
		4'd4: n_loc_oh_reg[217] = {11'd0, dist_reg[38], 4'd0};
		4'd5: n_loc_oh_reg[217] = {10'd0, dist_reg[38], 5'd0};
		4'd6: n_loc_oh_reg[217] = {9'd0, dist_reg[38], 6'd0};
		4'd7: n_loc_oh_reg[217] = {8'd0, dist_reg[38], 7'd0};
		4'd8: n_loc_oh_reg[217] = {7'd0, dist_reg[38], 8'd0};
		4'd9: n_loc_oh_reg[217] = {6'd0, dist_reg[38], 9'd0};
		4'd10: n_loc_oh_reg[217] = {5'd0, dist_reg[38], 10'd0};
		4'd11: n_loc_oh_reg[217] = {4'd0, dist_reg[38], 11'd0};
		4'd12: n_loc_oh_reg[217] = {3'd0, dist_reg[38], 12'd0};
		4'd13: n_loc_oh_reg[217] = {2'd0, dist_reg[38], 13'd0};
		4'd14: n_loc_oh_reg[217] = {1'd0, dist_reg[38], 14'd0};
		4'd15: n_loc_oh_reg[217] = {dist_reg[38], 15'd0};
	endcase
	case(loc_reg[218])
		4'd0: n_loc_oh_reg[218] = {15'd0, dist_reg[37]};
		4'd1: n_loc_oh_reg[218] = {14'd0, dist_reg[37], 1'd0};
		4'd2: n_loc_oh_reg[218] = {13'd0, dist_reg[37], 2'd0};
		4'd3: n_loc_oh_reg[218] = {12'd0, dist_reg[37], 3'd0};
		4'd4: n_loc_oh_reg[218] = {11'd0, dist_reg[37], 4'd0};
		4'd5: n_loc_oh_reg[218] = {10'd0, dist_reg[37], 5'd0};
		4'd6: n_loc_oh_reg[218] = {9'd0, dist_reg[37], 6'd0};
		4'd7: n_loc_oh_reg[218] = {8'd0, dist_reg[37], 7'd0};
		4'd8: n_loc_oh_reg[218] = {7'd0, dist_reg[37], 8'd0};
		4'd9: n_loc_oh_reg[218] = {6'd0, dist_reg[37], 9'd0};
		4'd10: n_loc_oh_reg[218] = {5'd0, dist_reg[37], 10'd0};
		4'd11: n_loc_oh_reg[218] = {4'd0, dist_reg[37], 11'd0};
		4'd12: n_loc_oh_reg[218] = {3'd0, dist_reg[37], 12'd0};
		4'd13: n_loc_oh_reg[218] = {2'd0, dist_reg[37], 13'd0};
		4'd14: n_loc_oh_reg[218] = {1'd0, dist_reg[37], 14'd0};
		4'd15: n_loc_oh_reg[218] = {dist_reg[37], 15'd0};
	endcase
	case(loc_reg[219])
		4'd0: n_loc_oh_reg[219] = {15'd0, dist_reg[36]};
		4'd1: n_loc_oh_reg[219] = {14'd0, dist_reg[36], 1'd0};
		4'd2: n_loc_oh_reg[219] = {13'd0, dist_reg[36], 2'd0};
		4'd3: n_loc_oh_reg[219] = {12'd0, dist_reg[36], 3'd0};
		4'd4: n_loc_oh_reg[219] = {11'd0, dist_reg[36], 4'd0};
		4'd5: n_loc_oh_reg[219] = {10'd0, dist_reg[36], 5'd0};
		4'd6: n_loc_oh_reg[219] = {9'd0, dist_reg[36], 6'd0};
		4'd7: n_loc_oh_reg[219] = {8'd0, dist_reg[36], 7'd0};
		4'd8: n_loc_oh_reg[219] = {7'd0, dist_reg[36], 8'd0};
		4'd9: n_loc_oh_reg[219] = {6'd0, dist_reg[36], 9'd0};
		4'd10: n_loc_oh_reg[219] = {5'd0, dist_reg[36], 10'd0};
		4'd11: n_loc_oh_reg[219] = {4'd0, dist_reg[36], 11'd0};
		4'd12: n_loc_oh_reg[219] = {3'd0, dist_reg[36], 12'd0};
		4'd13: n_loc_oh_reg[219] = {2'd0, dist_reg[36], 13'd0};
		4'd14: n_loc_oh_reg[219] = {1'd0, dist_reg[36], 14'd0};
		4'd15: n_loc_oh_reg[219] = {dist_reg[36], 15'd0};
	endcase
	case(loc_reg[220])
		4'd0: n_loc_oh_reg[220] = {15'd0, dist_reg[35]};
		4'd1: n_loc_oh_reg[220] = {14'd0, dist_reg[35], 1'd0};
		4'd2: n_loc_oh_reg[220] = {13'd0, dist_reg[35], 2'd0};
		4'd3: n_loc_oh_reg[220] = {12'd0, dist_reg[35], 3'd0};
		4'd4: n_loc_oh_reg[220] = {11'd0, dist_reg[35], 4'd0};
		4'd5: n_loc_oh_reg[220] = {10'd0, dist_reg[35], 5'd0};
		4'd6: n_loc_oh_reg[220] = {9'd0, dist_reg[35], 6'd0};
		4'd7: n_loc_oh_reg[220] = {8'd0, dist_reg[35], 7'd0};
		4'd8: n_loc_oh_reg[220] = {7'd0, dist_reg[35], 8'd0};
		4'd9: n_loc_oh_reg[220] = {6'd0, dist_reg[35], 9'd0};
		4'd10: n_loc_oh_reg[220] = {5'd0, dist_reg[35], 10'd0};
		4'd11: n_loc_oh_reg[220] = {4'd0, dist_reg[35], 11'd0};
		4'd12: n_loc_oh_reg[220] = {3'd0, dist_reg[35], 12'd0};
		4'd13: n_loc_oh_reg[220] = {2'd0, dist_reg[35], 13'd0};
		4'd14: n_loc_oh_reg[220] = {1'd0, dist_reg[35], 14'd0};
		4'd15: n_loc_oh_reg[220] = {dist_reg[35], 15'd0};
	endcase
	case(loc_reg[221])
		4'd0: n_loc_oh_reg[221] = {15'd0, dist_reg[34]};
		4'd1: n_loc_oh_reg[221] = {14'd0, dist_reg[34], 1'd0};
		4'd2: n_loc_oh_reg[221] = {13'd0, dist_reg[34], 2'd0};
		4'd3: n_loc_oh_reg[221] = {12'd0, dist_reg[34], 3'd0};
		4'd4: n_loc_oh_reg[221] = {11'd0, dist_reg[34], 4'd0};
		4'd5: n_loc_oh_reg[221] = {10'd0, dist_reg[34], 5'd0};
		4'd6: n_loc_oh_reg[221] = {9'd0, dist_reg[34], 6'd0};
		4'd7: n_loc_oh_reg[221] = {8'd0, dist_reg[34], 7'd0};
		4'd8: n_loc_oh_reg[221] = {7'd0, dist_reg[34], 8'd0};
		4'd9: n_loc_oh_reg[221] = {6'd0, dist_reg[34], 9'd0};
		4'd10: n_loc_oh_reg[221] = {5'd0, dist_reg[34], 10'd0};
		4'd11: n_loc_oh_reg[221] = {4'd0, dist_reg[34], 11'd0};
		4'd12: n_loc_oh_reg[221] = {3'd0, dist_reg[34], 12'd0};
		4'd13: n_loc_oh_reg[221] = {2'd0, dist_reg[34], 13'd0};
		4'd14: n_loc_oh_reg[221] = {1'd0, dist_reg[34], 14'd0};
		4'd15: n_loc_oh_reg[221] = {dist_reg[34], 15'd0};
	endcase
	case(loc_reg[222])
		4'd0: n_loc_oh_reg[222] = {15'd0, dist_reg[33]};
		4'd1: n_loc_oh_reg[222] = {14'd0, dist_reg[33], 1'd0};
		4'd2: n_loc_oh_reg[222] = {13'd0, dist_reg[33], 2'd0};
		4'd3: n_loc_oh_reg[222] = {12'd0, dist_reg[33], 3'd0};
		4'd4: n_loc_oh_reg[222] = {11'd0, dist_reg[33], 4'd0};
		4'd5: n_loc_oh_reg[222] = {10'd0, dist_reg[33], 5'd0};
		4'd6: n_loc_oh_reg[222] = {9'd0, dist_reg[33], 6'd0};
		4'd7: n_loc_oh_reg[222] = {8'd0, dist_reg[33], 7'd0};
		4'd8: n_loc_oh_reg[222] = {7'd0, dist_reg[33], 8'd0};
		4'd9: n_loc_oh_reg[222] = {6'd0, dist_reg[33], 9'd0};
		4'd10: n_loc_oh_reg[222] = {5'd0, dist_reg[33], 10'd0};
		4'd11: n_loc_oh_reg[222] = {4'd0, dist_reg[33], 11'd0};
		4'd12: n_loc_oh_reg[222] = {3'd0, dist_reg[33], 12'd0};
		4'd13: n_loc_oh_reg[222] = {2'd0, dist_reg[33], 13'd0};
		4'd14: n_loc_oh_reg[222] = {1'd0, dist_reg[33], 14'd0};
		4'd15: n_loc_oh_reg[222] = {dist_reg[33], 15'd0};
	endcase
	case(loc_reg[223])
		4'd0: n_loc_oh_reg[223] = {15'd0, dist_reg[32]};
		4'd1: n_loc_oh_reg[223] = {14'd0, dist_reg[32], 1'd0};
		4'd2: n_loc_oh_reg[223] = {13'd0, dist_reg[32], 2'd0};
		4'd3: n_loc_oh_reg[223] = {12'd0, dist_reg[32], 3'd0};
		4'd4: n_loc_oh_reg[223] = {11'd0, dist_reg[32], 4'd0};
		4'd5: n_loc_oh_reg[223] = {10'd0, dist_reg[32], 5'd0};
		4'd6: n_loc_oh_reg[223] = {9'd0, dist_reg[32], 6'd0};
		4'd7: n_loc_oh_reg[223] = {8'd0, dist_reg[32], 7'd0};
		4'd8: n_loc_oh_reg[223] = {7'd0, dist_reg[32], 8'd0};
		4'd9: n_loc_oh_reg[223] = {6'd0, dist_reg[32], 9'd0};
		4'd10: n_loc_oh_reg[223] = {5'd0, dist_reg[32], 10'd0};
		4'd11: n_loc_oh_reg[223] = {4'd0, dist_reg[32], 11'd0};
		4'd12: n_loc_oh_reg[223] = {3'd0, dist_reg[32], 12'd0};
		4'd13: n_loc_oh_reg[223] = {2'd0, dist_reg[32], 13'd0};
		4'd14: n_loc_oh_reg[223] = {1'd0, dist_reg[32], 14'd0};
		4'd15: n_loc_oh_reg[223] = {dist_reg[32], 15'd0};
	endcase
	case(loc_reg[224])
		4'd0: n_loc_oh_reg[224] = {15'd0, dist_reg[31]};
		4'd1: n_loc_oh_reg[224] = {14'd0, dist_reg[31], 1'd0};
		4'd2: n_loc_oh_reg[224] = {13'd0, dist_reg[31], 2'd0};
		4'd3: n_loc_oh_reg[224] = {12'd0, dist_reg[31], 3'd0};
		4'd4: n_loc_oh_reg[224] = {11'd0, dist_reg[31], 4'd0};
		4'd5: n_loc_oh_reg[224] = {10'd0, dist_reg[31], 5'd0};
		4'd6: n_loc_oh_reg[224] = {9'd0, dist_reg[31], 6'd0};
		4'd7: n_loc_oh_reg[224] = {8'd0, dist_reg[31], 7'd0};
		4'd8: n_loc_oh_reg[224] = {7'd0, dist_reg[31], 8'd0};
		4'd9: n_loc_oh_reg[224] = {6'd0, dist_reg[31], 9'd0};
		4'd10: n_loc_oh_reg[224] = {5'd0, dist_reg[31], 10'd0};
		4'd11: n_loc_oh_reg[224] = {4'd0, dist_reg[31], 11'd0};
		4'd12: n_loc_oh_reg[224] = {3'd0, dist_reg[31], 12'd0};
		4'd13: n_loc_oh_reg[224] = {2'd0, dist_reg[31], 13'd0};
		4'd14: n_loc_oh_reg[224] = {1'd0, dist_reg[31], 14'd0};
		4'd15: n_loc_oh_reg[224] = {dist_reg[31], 15'd0};
	endcase
	case(loc_reg[225])
		4'd0: n_loc_oh_reg[225] = {15'd0, dist_reg[30]};
		4'd1: n_loc_oh_reg[225] = {14'd0, dist_reg[30], 1'd0};
		4'd2: n_loc_oh_reg[225] = {13'd0, dist_reg[30], 2'd0};
		4'd3: n_loc_oh_reg[225] = {12'd0, dist_reg[30], 3'd0};
		4'd4: n_loc_oh_reg[225] = {11'd0, dist_reg[30], 4'd0};
		4'd5: n_loc_oh_reg[225] = {10'd0, dist_reg[30], 5'd0};
		4'd6: n_loc_oh_reg[225] = {9'd0, dist_reg[30], 6'd0};
		4'd7: n_loc_oh_reg[225] = {8'd0, dist_reg[30], 7'd0};
		4'd8: n_loc_oh_reg[225] = {7'd0, dist_reg[30], 8'd0};
		4'd9: n_loc_oh_reg[225] = {6'd0, dist_reg[30], 9'd0};
		4'd10: n_loc_oh_reg[225] = {5'd0, dist_reg[30], 10'd0};
		4'd11: n_loc_oh_reg[225] = {4'd0, dist_reg[30], 11'd0};
		4'd12: n_loc_oh_reg[225] = {3'd0, dist_reg[30], 12'd0};
		4'd13: n_loc_oh_reg[225] = {2'd0, dist_reg[30], 13'd0};
		4'd14: n_loc_oh_reg[225] = {1'd0, dist_reg[30], 14'd0};
		4'd15: n_loc_oh_reg[225] = {dist_reg[30], 15'd0};
	endcase
	case(loc_reg[226])
		4'd0: n_loc_oh_reg[226] = {15'd0, dist_reg[29]};
		4'd1: n_loc_oh_reg[226] = {14'd0, dist_reg[29], 1'd0};
		4'd2: n_loc_oh_reg[226] = {13'd0, dist_reg[29], 2'd0};
		4'd3: n_loc_oh_reg[226] = {12'd0, dist_reg[29], 3'd0};
		4'd4: n_loc_oh_reg[226] = {11'd0, dist_reg[29], 4'd0};
		4'd5: n_loc_oh_reg[226] = {10'd0, dist_reg[29], 5'd0};
		4'd6: n_loc_oh_reg[226] = {9'd0, dist_reg[29], 6'd0};
		4'd7: n_loc_oh_reg[226] = {8'd0, dist_reg[29], 7'd0};
		4'd8: n_loc_oh_reg[226] = {7'd0, dist_reg[29], 8'd0};
		4'd9: n_loc_oh_reg[226] = {6'd0, dist_reg[29], 9'd0};
		4'd10: n_loc_oh_reg[226] = {5'd0, dist_reg[29], 10'd0};
		4'd11: n_loc_oh_reg[226] = {4'd0, dist_reg[29], 11'd0};
		4'd12: n_loc_oh_reg[226] = {3'd0, dist_reg[29], 12'd0};
		4'd13: n_loc_oh_reg[226] = {2'd0, dist_reg[29], 13'd0};
		4'd14: n_loc_oh_reg[226] = {1'd0, dist_reg[29], 14'd0};
		4'd15: n_loc_oh_reg[226] = {dist_reg[29], 15'd0};
	endcase
	case(loc_reg[227])
		4'd0: n_loc_oh_reg[227] = {15'd0, dist_reg[28]};
		4'd1: n_loc_oh_reg[227] = {14'd0, dist_reg[28], 1'd0};
		4'd2: n_loc_oh_reg[227] = {13'd0, dist_reg[28], 2'd0};
		4'd3: n_loc_oh_reg[227] = {12'd0, dist_reg[28], 3'd0};
		4'd4: n_loc_oh_reg[227] = {11'd0, dist_reg[28], 4'd0};
		4'd5: n_loc_oh_reg[227] = {10'd0, dist_reg[28], 5'd0};
		4'd6: n_loc_oh_reg[227] = {9'd0, dist_reg[28], 6'd0};
		4'd7: n_loc_oh_reg[227] = {8'd0, dist_reg[28], 7'd0};
		4'd8: n_loc_oh_reg[227] = {7'd0, dist_reg[28], 8'd0};
		4'd9: n_loc_oh_reg[227] = {6'd0, dist_reg[28], 9'd0};
		4'd10: n_loc_oh_reg[227] = {5'd0, dist_reg[28], 10'd0};
		4'd11: n_loc_oh_reg[227] = {4'd0, dist_reg[28], 11'd0};
		4'd12: n_loc_oh_reg[227] = {3'd0, dist_reg[28], 12'd0};
		4'd13: n_loc_oh_reg[227] = {2'd0, dist_reg[28], 13'd0};
		4'd14: n_loc_oh_reg[227] = {1'd0, dist_reg[28], 14'd0};
		4'd15: n_loc_oh_reg[227] = {dist_reg[28], 15'd0};
	endcase
	case(loc_reg[228])
		4'd0: n_loc_oh_reg[228] = {15'd0, dist_reg[27]};
		4'd1: n_loc_oh_reg[228] = {14'd0, dist_reg[27], 1'd0};
		4'd2: n_loc_oh_reg[228] = {13'd0, dist_reg[27], 2'd0};
		4'd3: n_loc_oh_reg[228] = {12'd0, dist_reg[27], 3'd0};
		4'd4: n_loc_oh_reg[228] = {11'd0, dist_reg[27], 4'd0};
		4'd5: n_loc_oh_reg[228] = {10'd0, dist_reg[27], 5'd0};
		4'd6: n_loc_oh_reg[228] = {9'd0, dist_reg[27], 6'd0};
		4'd7: n_loc_oh_reg[228] = {8'd0, dist_reg[27], 7'd0};
		4'd8: n_loc_oh_reg[228] = {7'd0, dist_reg[27], 8'd0};
		4'd9: n_loc_oh_reg[228] = {6'd0, dist_reg[27], 9'd0};
		4'd10: n_loc_oh_reg[228] = {5'd0, dist_reg[27], 10'd0};
		4'd11: n_loc_oh_reg[228] = {4'd0, dist_reg[27], 11'd0};
		4'd12: n_loc_oh_reg[228] = {3'd0, dist_reg[27], 12'd0};
		4'd13: n_loc_oh_reg[228] = {2'd0, dist_reg[27], 13'd0};
		4'd14: n_loc_oh_reg[228] = {1'd0, dist_reg[27], 14'd0};
		4'd15: n_loc_oh_reg[228] = {dist_reg[27], 15'd0};
	endcase
	case(loc_reg[229])
		4'd0: n_loc_oh_reg[229] = {15'd0, dist_reg[26]};
		4'd1: n_loc_oh_reg[229] = {14'd0, dist_reg[26], 1'd0};
		4'd2: n_loc_oh_reg[229] = {13'd0, dist_reg[26], 2'd0};
		4'd3: n_loc_oh_reg[229] = {12'd0, dist_reg[26], 3'd0};
		4'd4: n_loc_oh_reg[229] = {11'd0, dist_reg[26], 4'd0};
		4'd5: n_loc_oh_reg[229] = {10'd0, dist_reg[26], 5'd0};
		4'd6: n_loc_oh_reg[229] = {9'd0, dist_reg[26], 6'd0};
		4'd7: n_loc_oh_reg[229] = {8'd0, dist_reg[26], 7'd0};
		4'd8: n_loc_oh_reg[229] = {7'd0, dist_reg[26], 8'd0};
		4'd9: n_loc_oh_reg[229] = {6'd0, dist_reg[26], 9'd0};
		4'd10: n_loc_oh_reg[229] = {5'd0, dist_reg[26], 10'd0};
		4'd11: n_loc_oh_reg[229] = {4'd0, dist_reg[26], 11'd0};
		4'd12: n_loc_oh_reg[229] = {3'd0, dist_reg[26], 12'd0};
		4'd13: n_loc_oh_reg[229] = {2'd0, dist_reg[26], 13'd0};
		4'd14: n_loc_oh_reg[229] = {1'd0, dist_reg[26], 14'd0};
		4'd15: n_loc_oh_reg[229] = {dist_reg[26], 15'd0};
	endcase
	case(loc_reg[230])
		4'd0: n_loc_oh_reg[230] = {15'd0, dist_reg[25]};
		4'd1: n_loc_oh_reg[230] = {14'd0, dist_reg[25], 1'd0};
		4'd2: n_loc_oh_reg[230] = {13'd0, dist_reg[25], 2'd0};
		4'd3: n_loc_oh_reg[230] = {12'd0, dist_reg[25], 3'd0};
		4'd4: n_loc_oh_reg[230] = {11'd0, dist_reg[25], 4'd0};
		4'd5: n_loc_oh_reg[230] = {10'd0, dist_reg[25], 5'd0};
		4'd6: n_loc_oh_reg[230] = {9'd0, dist_reg[25], 6'd0};
		4'd7: n_loc_oh_reg[230] = {8'd0, dist_reg[25], 7'd0};
		4'd8: n_loc_oh_reg[230] = {7'd0, dist_reg[25], 8'd0};
		4'd9: n_loc_oh_reg[230] = {6'd0, dist_reg[25], 9'd0};
		4'd10: n_loc_oh_reg[230] = {5'd0, dist_reg[25], 10'd0};
		4'd11: n_loc_oh_reg[230] = {4'd0, dist_reg[25], 11'd0};
		4'd12: n_loc_oh_reg[230] = {3'd0, dist_reg[25], 12'd0};
		4'd13: n_loc_oh_reg[230] = {2'd0, dist_reg[25], 13'd0};
		4'd14: n_loc_oh_reg[230] = {1'd0, dist_reg[25], 14'd0};
		4'd15: n_loc_oh_reg[230] = {dist_reg[25], 15'd0};
	endcase
	case(loc_reg[231])
		4'd0: n_loc_oh_reg[231] = {15'd0, dist_reg[24]};
		4'd1: n_loc_oh_reg[231] = {14'd0, dist_reg[24], 1'd0};
		4'd2: n_loc_oh_reg[231] = {13'd0, dist_reg[24], 2'd0};
		4'd3: n_loc_oh_reg[231] = {12'd0, dist_reg[24], 3'd0};
		4'd4: n_loc_oh_reg[231] = {11'd0, dist_reg[24], 4'd0};
		4'd5: n_loc_oh_reg[231] = {10'd0, dist_reg[24], 5'd0};
		4'd6: n_loc_oh_reg[231] = {9'd0, dist_reg[24], 6'd0};
		4'd7: n_loc_oh_reg[231] = {8'd0, dist_reg[24], 7'd0};
		4'd8: n_loc_oh_reg[231] = {7'd0, dist_reg[24], 8'd0};
		4'd9: n_loc_oh_reg[231] = {6'd0, dist_reg[24], 9'd0};
		4'd10: n_loc_oh_reg[231] = {5'd0, dist_reg[24], 10'd0};
		4'd11: n_loc_oh_reg[231] = {4'd0, dist_reg[24], 11'd0};
		4'd12: n_loc_oh_reg[231] = {3'd0, dist_reg[24], 12'd0};
		4'd13: n_loc_oh_reg[231] = {2'd0, dist_reg[24], 13'd0};
		4'd14: n_loc_oh_reg[231] = {1'd0, dist_reg[24], 14'd0};
		4'd15: n_loc_oh_reg[231] = {dist_reg[24], 15'd0};
	endcase
	case(loc_reg[232])
		4'd0: n_loc_oh_reg[232] = {15'd0, dist_reg[23]};
		4'd1: n_loc_oh_reg[232] = {14'd0, dist_reg[23], 1'd0};
		4'd2: n_loc_oh_reg[232] = {13'd0, dist_reg[23], 2'd0};
		4'd3: n_loc_oh_reg[232] = {12'd0, dist_reg[23], 3'd0};
		4'd4: n_loc_oh_reg[232] = {11'd0, dist_reg[23], 4'd0};
		4'd5: n_loc_oh_reg[232] = {10'd0, dist_reg[23], 5'd0};
		4'd6: n_loc_oh_reg[232] = {9'd0, dist_reg[23], 6'd0};
		4'd7: n_loc_oh_reg[232] = {8'd0, dist_reg[23], 7'd0};
		4'd8: n_loc_oh_reg[232] = {7'd0, dist_reg[23], 8'd0};
		4'd9: n_loc_oh_reg[232] = {6'd0, dist_reg[23], 9'd0};
		4'd10: n_loc_oh_reg[232] = {5'd0, dist_reg[23], 10'd0};
		4'd11: n_loc_oh_reg[232] = {4'd0, dist_reg[23], 11'd0};
		4'd12: n_loc_oh_reg[232] = {3'd0, dist_reg[23], 12'd0};
		4'd13: n_loc_oh_reg[232] = {2'd0, dist_reg[23], 13'd0};
		4'd14: n_loc_oh_reg[232] = {1'd0, dist_reg[23], 14'd0};
		4'd15: n_loc_oh_reg[232] = {dist_reg[23], 15'd0};
	endcase
	case(loc_reg[233])
		4'd0: n_loc_oh_reg[233] = {15'd0, dist_reg[22]};
		4'd1: n_loc_oh_reg[233] = {14'd0, dist_reg[22], 1'd0};
		4'd2: n_loc_oh_reg[233] = {13'd0, dist_reg[22], 2'd0};
		4'd3: n_loc_oh_reg[233] = {12'd0, dist_reg[22], 3'd0};
		4'd4: n_loc_oh_reg[233] = {11'd0, dist_reg[22], 4'd0};
		4'd5: n_loc_oh_reg[233] = {10'd0, dist_reg[22], 5'd0};
		4'd6: n_loc_oh_reg[233] = {9'd0, dist_reg[22], 6'd0};
		4'd7: n_loc_oh_reg[233] = {8'd0, dist_reg[22], 7'd0};
		4'd8: n_loc_oh_reg[233] = {7'd0, dist_reg[22], 8'd0};
		4'd9: n_loc_oh_reg[233] = {6'd0, dist_reg[22], 9'd0};
		4'd10: n_loc_oh_reg[233] = {5'd0, dist_reg[22], 10'd0};
		4'd11: n_loc_oh_reg[233] = {4'd0, dist_reg[22], 11'd0};
		4'd12: n_loc_oh_reg[233] = {3'd0, dist_reg[22], 12'd0};
		4'd13: n_loc_oh_reg[233] = {2'd0, dist_reg[22], 13'd0};
		4'd14: n_loc_oh_reg[233] = {1'd0, dist_reg[22], 14'd0};
		4'd15: n_loc_oh_reg[233] = {dist_reg[22], 15'd0};
	endcase
	case(loc_reg[234])
		4'd0: n_loc_oh_reg[234] = {15'd0, dist_reg[21]};
		4'd1: n_loc_oh_reg[234] = {14'd0, dist_reg[21], 1'd0};
		4'd2: n_loc_oh_reg[234] = {13'd0, dist_reg[21], 2'd0};
		4'd3: n_loc_oh_reg[234] = {12'd0, dist_reg[21], 3'd0};
		4'd4: n_loc_oh_reg[234] = {11'd0, dist_reg[21], 4'd0};
		4'd5: n_loc_oh_reg[234] = {10'd0, dist_reg[21], 5'd0};
		4'd6: n_loc_oh_reg[234] = {9'd0, dist_reg[21], 6'd0};
		4'd7: n_loc_oh_reg[234] = {8'd0, dist_reg[21], 7'd0};
		4'd8: n_loc_oh_reg[234] = {7'd0, dist_reg[21], 8'd0};
		4'd9: n_loc_oh_reg[234] = {6'd0, dist_reg[21], 9'd0};
		4'd10: n_loc_oh_reg[234] = {5'd0, dist_reg[21], 10'd0};
		4'd11: n_loc_oh_reg[234] = {4'd0, dist_reg[21], 11'd0};
		4'd12: n_loc_oh_reg[234] = {3'd0, dist_reg[21], 12'd0};
		4'd13: n_loc_oh_reg[234] = {2'd0, dist_reg[21], 13'd0};
		4'd14: n_loc_oh_reg[234] = {1'd0, dist_reg[21], 14'd0};
		4'd15: n_loc_oh_reg[234] = {dist_reg[21], 15'd0};
	endcase
	case(loc_reg[235])
		4'd0: n_loc_oh_reg[235] = {15'd0, dist_reg[20]};
		4'd1: n_loc_oh_reg[235] = {14'd0, dist_reg[20], 1'd0};
		4'd2: n_loc_oh_reg[235] = {13'd0, dist_reg[20], 2'd0};
		4'd3: n_loc_oh_reg[235] = {12'd0, dist_reg[20], 3'd0};
		4'd4: n_loc_oh_reg[235] = {11'd0, dist_reg[20], 4'd0};
		4'd5: n_loc_oh_reg[235] = {10'd0, dist_reg[20], 5'd0};
		4'd6: n_loc_oh_reg[235] = {9'd0, dist_reg[20], 6'd0};
		4'd7: n_loc_oh_reg[235] = {8'd0, dist_reg[20], 7'd0};
		4'd8: n_loc_oh_reg[235] = {7'd0, dist_reg[20], 8'd0};
		4'd9: n_loc_oh_reg[235] = {6'd0, dist_reg[20], 9'd0};
		4'd10: n_loc_oh_reg[235] = {5'd0, dist_reg[20], 10'd0};
		4'd11: n_loc_oh_reg[235] = {4'd0, dist_reg[20], 11'd0};
		4'd12: n_loc_oh_reg[235] = {3'd0, dist_reg[20], 12'd0};
		4'd13: n_loc_oh_reg[235] = {2'd0, dist_reg[20], 13'd0};
		4'd14: n_loc_oh_reg[235] = {1'd0, dist_reg[20], 14'd0};
		4'd15: n_loc_oh_reg[235] = {dist_reg[20], 15'd0};
	endcase
	case(loc_reg[236])
		4'd0: n_loc_oh_reg[236] = {15'd0, dist_reg[19]};
		4'd1: n_loc_oh_reg[236] = {14'd0, dist_reg[19], 1'd0};
		4'd2: n_loc_oh_reg[236] = {13'd0, dist_reg[19], 2'd0};
		4'd3: n_loc_oh_reg[236] = {12'd0, dist_reg[19], 3'd0};
		4'd4: n_loc_oh_reg[236] = {11'd0, dist_reg[19], 4'd0};
		4'd5: n_loc_oh_reg[236] = {10'd0, dist_reg[19], 5'd0};
		4'd6: n_loc_oh_reg[236] = {9'd0, dist_reg[19], 6'd0};
		4'd7: n_loc_oh_reg[236] = {8'd0, dist_reg[19], 7'd0};
		4'd8: n_loc_oh_reg[236] = {7'd0, dist_reg[19], 8'd0};
		4'd9: n_loc_oh_reg[236] = {6'd0, dist_reg[19], 9'd0};
		4'd10: n_loc_oh_reg[236] = {5'd0, dist_reg[19], 10'd0};
		4'd11: n_loc_oh_reg[236] = {4'd0, dist_reg[19], 11'd0};
		4'd12: n_loc_oh_reg[236] = {3'd0, dist_reg[19], 12'd0};
		4'd13: n_loc_oh_reg[236] = {2'd0, dist_reg[19], 13'd0};
		4'd14: n_loc_oh_reg[236] = {1'd0, dist_reg[19], 14'd0};
		4'd15: n_loc_oh_reg[236] = {dist_reg[19], 15'd0};
	endcase
	case(loc_reg[237])
		4'd0: n_loc_oh_reg[237] = {15'd0, dist_reg[18]};
		4'd1: n_loc_oh_reg[237] = {14'd0, dist_reg[18], 1'd0};
		4'd2: n_loc_oh_reg[237] = {13'd0, dist_reg[18], 2'd0};
		4'd3: n_loc_oh_reg[237] = {12'd0, dist_reg[18], 3'd0};
		4'd4: n_loc_oh_reg[237] = {11'd0, dist_reg[18], 4'd0};
		4'd5: n_loc_oh_reg[237] = {10'd0, dist_reg[18], 5'd0};
		4'd6: n_loc_oh_reg[237] = {9'd0, dist_reg[18], 6'd0};
		4'd7: n_loc_oh_reg[237] = {8'd0, dist_reg[18], 7'd0};
		4'd8: n_loc_oh_reg[237] = {7'd0, dist_reg[18], 8'd0};
		4'd9: n_loc_oh_reg[237] = {6'd0, dist_reg[18], 9'd0};
		4'd10: n_loc_oh_reg[237] = {5'd0, dist_reg[18], 10'd0};
		4'd11: n_loc_oh_reg[237] = {4'd0, dist_reg[18], 11'd0};
		4'd12: n_loc_oh_reg[237] = {3'd0, dist_reg[18], 12'd0};
		4'd13: n_loc_oh_reg[237] = {2'd0, dist_reg[18], 13'd0};
		4'd14: n_loc_oh_reg[237] = {1'd0, dist_reg[18], 14'd0};
		4'd15: n_loc_oh_reg[237] = {dist_reg[18], 15'd0};
	endcase
	case(loc_reg[238])
		4'd0: n_loc_oh_reg[238] = {15'd0, dist_reg[17]};
		4'd1: n_loc_oh_reg[238] = {14'd0, dist_reg[17], 1'd0};
		4'd2: n_loc_oh_reg[238] = {13'd0, dist_reg[17], 2'd0};
		4'd3: n_loc_oh_reg[238] = {12'd0, dist_reg[17], 3'd0};
		4'd4: n_loc_oh_reg[238] = {11'd0, dist_reg[17], 4'd0};
		4'd5: n_loc_oh_reg[238] = {10'd0, dist_reg[17], 5'd0};
		4'd6: n_loc_oh_reg[238] = {9'd0, dist_reg[17], 6'd0};
		4'd7: n_loc_oh_reg[238] = {8'd0, dist_reg[17], 7'd0};
		4'd8: n_loc_oh_reg[238] = {7'd0, dist_reg[17], 8'd0};
		4'd9: n_loc_oh_reg[238] = {6'd0, dist_reg[17], 9'd0};
		4'd10: n_loc_oh_reg[238] = {5'd0, dist_reg[17], 10'd0};
		4'd11: n_loc_oh_reg[238] = {4'd0, dist_reg[17], 11'd0};
		4'd12: n_loc_oh_reg[238] = {3'd0, dist_reg[17], 12'd0};
		4'd13: n_loc_oh_reg[238] = {2'd0, dist_reg[17], 13'd0};
		4'd14: n_loc_oh_reg[238] = {1'd0, dist_reg[17], 14'd0};
		4'd15: n_loc_oh_reg[238] = {dist_reg[17], 15'd0};
	endcase
	case(loc_reg[239])
		4'd0: n_loc_oh_reg[239] = {15'd0, dist_reg[16]};
		4'd1: n_loc_oh_reg[239] = {14'd0, dist_reg[16], 1'd0};
		4'd2: n_loc_oh_reg[239] = {13'd0, dist_reg[16], 2'd0};
		4'd3: n_loc_oh_reg[239] = {12'd0, dist_reg[16], 3'd0};
		4'd4: n_loc_oh_reg[239] = {11'd0, dist_reg[16], 4'd0};
		4'd5: n_loc_oh_reg[239] = {10'd0, dist_reg[16], 5'd0};
		4'd6: n_loc_oh_reg[239] = {9'd0, dist_reg[16], 6'd0};
		4'd7: n_loc_oh_reg[239] = {8'd0, dist_reg[16], 7'd0};
		4'd8: n_loc_oh_reg[239] = {7'd0, dist_reg[16], 8'd0};
		4'd9: n_loc_oh_reg[239] = {6'd0, dist_reg[16], 9'd0};
		4'd10: n_loc_oh_reg[239] = {5'd0, dist_reg[16], 10'd0};
		4'd11: n_loc_oh_reg[239] = {4'd0, dist_reg[16], 11'd0};
		4'd12: n_loc_oh_reg[239] = {3'd0, dist_reg[16], 12'd0};
		4'd13: n_loc_oh_reg[239] = {2'd0, dist_reg[16], 13'd0};
		4'd14: n_loc_oh_reg[239] = {1'd0, dist_reg[16], 14'd0};
		4'd15: n_loc_oh_reg[239] = {dist_reg[16], 15'd0};
	endcase
	case(loc_reg[240])
		4'd0: n_loc_oh_reg[240] = {15'd0, dist_reg[15]};
		4'd1: n_loc_oh_reg[240] = {14'd0, dist_reg[15], 1'd0};
		4'd2: n_loc_oh_reg[240] = {13'd0, dist_reg[15], 2'd0};
		4'd3: n_loc_oh_reg[240] = {12'd0, dist_reg[15], 3'd0};
		4'd4: n_loc_oh_reg[240] = {11'd0, dist_reg[15], 4'd0};
		4'd5: n_loc_oh_reg[240] = {10'd0, dist_reg[15], 5'd0};
		4'd6: n_loc_oh_reg[240] = {9'd0, dist_reg[15], 6'd0};
		4'd7: n_loc_oh_reg[240] = {8'd0, dist_reg[15], 7'd0};
		4'd8: n_loc_oh_reg[240] = {7'd0, dist_reg[15], 8'd0};
		4'd9: n_loc_oh_reg[240] = {6'd0, dist_reg[15], 9'd0};
		4'd10: n_loc_oh_reg[240] = {5'd0, dist_reg[15], 10'd0};
		4'd11: n_loc_oh_reg[240] = {4'd0, dist_reg[15], 11'd0};
		4'd12: n_loc_oh_reg[240] = {3'd0, dist_reg[15], 12'd0};
		4'd13: n_loc_oh_reg[240] = {2'd0, dist_reg[15], 13'd0};
		4'd14: n_loc_oh_reg[240] = {1'd0, dist_reg[15], 14'd0};
		4'd15: n_loc_oh_reg[240] = {dist_reg[15], 15'd0};
	endcase
	case(loc_reg[241])
		4'd0: n_loc_oh_reg[241] = {15'd0, dist_reg[14]};
		4'd1: n_loc_oh_reg[241] = {14'd0, dist_reg[14], 1'd0};
		4'd2: n_loc_oh_reg[241] = {13'd0, dist_reg[14], 2'd0};
		4'd3: n_loc_oh_reg[241] = {12'd0, dist_reg[14], 3'd0};
		4'd4: n_loc_oh_reg[241] = {11'd0, dist_reg[14], 4'd0};
		4'd5: n_loc_oh_reg[241] = {10'd0, dist_reg[14], 5'd0};
		4'd6: n_loc_oh_reg[241] = {9'd0, dist_reg[14], 6'd0};
		4'd7: n_loc_oh_reg[241] = {8'd0, dist_reg[14], 7'd0};
		4'd8: n_loc_oh_reg[241] = {7'd0, dist_reg[14], 8'd0};
		4'd9: n_loc_oh_reg[241] = {6'd0, dist_reg[14], 9'd0};
		4'd10: n_loc_oh_reg[241] = {5'd0, dist_reg[14], 10'd0};
		4'd11: n_loc_oh_reg[241] = {4'd0, dist_reg[14], 11'd0};
		4'd12: n_loc_oh_reg[241] = {3'd0, dist_reg[14], 12'd0};
		4'd13: n_loc_oh_reg[241] = {2'd0, dist_reg[14], 13'd0};
		4'd14: n_loc_oh_reg[241] = {1'd0, dist_reg[14], 14'd0};
		4'd15: n_loc_oh_reg[241] = {dist_reg[14], 15'd0};
	endcase
	case(loc_reg[242])
		4'd0: n_loc_oh_reg[242] = {15'd0, dist_reg[13]};
		4'd1: n_loc_oh_reg[242] = {14'd0, dist_reg[13], 1'd0};
		4'd2: n_loc_oh_reg[242] = {13'd0, dist_reg[13], 2'd0};
		4'd3: n_loc_oh_reg[242] = {12'd0, dist_reg[13], 3'd0};
		4'd4: n_loc_oh_reg[242] = {11'd0, dist_reg[13], 4'd0};
		4'd5: n_loc_oh_reg[242] = {10'd0, dist_reg[13], 5'd0};
		4'd6: n_loc_oh_reg[242] = {9'd0, dist_reg[13], 6'd0};
		4'd7: n_loc_oh_reg[242] = {8'd0, dist_reg[13], 7'd0};
		4'd8: n_loc_oh_reg[242] = {7'd0, dist_reg[13], 8'd0};
		4'd9: n_loc_oh_reg[242] = {6'd0, dist_reg[13], 9'd0};
		4'd10: n_loc_oh_reg[242] = {5'd0, dist_reg[13], 10'd0};
		4'd11: n_loc_oh_reg[242] = {4'd0, dist_reg[13], 11'd0};
		4'd12: n_loc_oh_reg[242] = {3'd0, dist_reg[13], 12'd0};
		4'd13: n_loc_oh_reg[242] = {2'd0, dist_reg[13], 13'd0};
		4'd14: n_loc_oh_reg[242] = {1'd0, dist_reg[13], 14'd0};
		4'd15: n_loc_oh_reg[242] = {dist_reg[13], 15'd0};
	endcase
	case(loc_reg[243])
		4'd0: n_loc_oh_reg[243] = {15'd0, dist_reg[12]};
		4'd1: n_loc_oh_reg[243] = {14'd0, dist_reg[12], 1'd0};
		4'd2: n_loc_oh_reg[243] = {13'd0, dist_reg[12], 2'd0};
		4'd3: n_loc_oh_reg[243] = {12'd0, dist_reg[12], 3'd0};
		4'd4: n_loc_oh_reg[243] = {11'd0, dist_reg[12], 4'd0};
		4'd5: n_loc_oh_reg[243] = {10'd0, dist_reg[12], 5'd0};
		4'd6: n_loc_oh_reg[243] = {9'd0, dist_reg[12], 6'd0};
		4'd7: n_loc_oh_reg[243] = {8'd0, dist_reg[12], 7'd0};
		4'd8: n_loc_oh_reg[243] = {7'd0, dist_reg[12], 8'd0};
		4'd9: n_loc_oh_reg[243] = {6'd0, dist_reg[12], 9'd0};
		4'd10: n_loc_oh_reg[243] = {5'd0, dist_reg[12], 10'd0};
		4'd11: n_loc_oh_reg[243] = {4'd0, dist_reg[12], 11'd0};
		4'd12: n_loc_oh_reg[243] = {3'd0, dist_reg[12], 12'd0};
		4'd13: n_loc_oh_reg[243] = {2'd0, dist_reg[12], 13'd0};
		4'd14: n_loc_oh_reg[243] = {1'd0, dist_reg[12], 14'd0};
		4'd15: n_loc_oh_reg[243] = {dist_reg[12], 15'd0};
	endcase
	case(loc_reg[244])
		4'd0: n_loc_oh_reg[244] = {15'd0, dist_reg[11]};
		4'd1: n_loc_oh_reg[244] = {14'd0, dist_reg[11], 1'd0};
		4'd2: n_loc_oh_reg[244] = {13'd0, dist_reg[11], 2'd0};
		4'd3: n_loc_oh_reg[244] = {12'd0, dist_reg[11], 3'd0};
		4'd4: n_loc_oh_reg[244] = {11'd0, dist_reg[11], 4'd0};
		4'd5: n_loc_oh_reg[244] = {10'd0, dist_reg[11], 5'd0};
		4'd6: n_loc_oh_reg[244] = {9'd0, dist_reg[11], 6'd0};
		4'd7: n_loc_oh_reg[244] = {8'd0, dist_reg[11], 7'd0};
		4'd8: n_loc_oh_reg[244] = {7'd0, dist_reg[11], 8'd0};
		4'd9: n_loc_oh_reg[244] = {6'd0, dist_reg[11], 9'd0};
		4'd10: n_loc_oh_reg[244] = {5'd0, dist_reg[11], 10'd0};
		4'd11: n_loc_oh_reg[244] = {4'd0, dist_reg[11], 11'd0};
		4'd12: n_loc_oh_reg[244] = {3'd0, dist_reg[11], 12'd0};
		4'd13: n_loc_oh_reg[244] = {2'd0, dist_reg[11], 13'd0};
		4'd14: n_loc_oh_reg[244] = {1'd0, dist_reg[11], 14'd0};
		4'd15: n_loc_oh_reg[244] = {dist_reg[11], 15'd0};
	endcase
	case(loc_reg[245])
		4'd0: n_loc_oh_reg[245] = {15'd0, dist_reg[10]};
		4'd1: n_loc_oh_reg[245] = {14'd0, dist_reg[10], 1'd0};
		4'd2: n_loc_oh_reg[245] = {13'd0, dist_reg[10], 2'd0};
		4'd3: n_loc_oh_reg[245] = {12'd0, dist_reg[10], 3'd0};
		4'd4: n_loc_oh_reg[245] = {11'd0, dist_reg[10], 4'd0};
		4'd5: n_loc_oh_reg[245] = {10'd0, dist_reg[10], 5'd0};
		4'd6: n_loc_oh_reg[245] = {9'd0, dist_reg[10], 6'd0};
		4'd7: n_loc_oh_reg[245] = {8'd0, dist_reg[10], 7'd0};
		4'd8: n_loc_oh_reg[245] = {7'd0, dist_reg[10], 8'd0};
		4'd9: n_loc_oh_reg[245] = {6'd0, dist_reg[10], 9'd0};
		4'd10: n_loc_oh_reg[245] = {5'd0, dist_reg[10], 10'd0};
		4'd11: n_loc_oh_reg[245] = {4'd0, dist_reg[10], 11'd0};
		4'd12: n_loc_oh_reg[245] = {3'd0, dist_reg[10], 12'd0};
		4'd13: n_loc_oh_reg[245] = {2'd0, dist_reg[10], 13'd0};
		4'd14: n_loc_oh_reg[245] = {1'd0, dist_reg[10], 14'd0};
		4'd15: n_loc_oh_reg[245] = {dist_reg[10], 15'd0};
	endcase
	case(loc_reg[246])
		4'd0: n_loc_oh_reg[246] = {15'd0, dist_reg[9]};
		4'd1: n_loc_oh_reg[246] = {14'd0, dist_reg[9], 1'd0};
		4'd2: n_loc_oh_reg[246] = {13'd0, dist_reg[9], 2'd0};
		4'd3: n_loc_oh_reg[246] = {12'd0, dist_reg[9], 3'd0};
		4'd4: n_loc_oh_reg[246] = {11'd0, dist_reg[9], 4'd0};
		4'd5: n_loc_oh_reg[246] = {10'd0, dist_reg[9], 5'd0};
		4'd6: n_loc_oh_reg[246] = {9'd0, dist_reg[9], 6'd0};
		4'd7: n_loc_oh_reg[246] = {8'd0, dist_reg[9], 7'd0};
		4'd8: n_loc_oh_reg[246] = {7'd0, dist_reg[9], 8'd0};
		4'd9: n_loc_oh_reg[246] = {6'd0, dist_reg[9], 9'd0};
		4'd10: n_loc_oh_reg[246] = {5'd0, dist_reg[9], 10'd0};
		4'd11: n_loc_oh_reg[246] = {4'd0, dist_reg[9], 11'd0};
		4'd12: n_loc_oh_reg[246] = {3'd0, dist_reg[9], 12'd0};
		4'd13: n_loc_oh_reg[246] = {2'd0, dist_reg[9], 13'd0};
		4'd14: n_loc_oh_reg[246] = {1'd0, dist_reg[9], 14'd0};
		4'd15: n_loc_oh_reg[246] = {dist_reg[9], 15'd0};
	endcase
	case(loc_reg[247])
		4'd0: n_loc_oh_reg[247] = {15'd0, dist_reg[8]};
		4'd1: n_loc_oh_reg[247] = {14'd0, dist_reg[8], 1'd0};
		4'd2: n_loc_oh_reg[247] = {13'd0, dist_reg[8], 2'd0};
		4'd3: n_loc_oh_reg[247] = {12'd0, dist_reg[8], 3'd0};
		4'd4: n_loc_oh_reg[247] = {11'd0, dist_reg[8], 4'd0};
		4'd5: n_loc_oh_reg[247] = {10'd0, dist_reg[8], 5'd0};
		4'd6: n_loc_oh_reg[247] = {9'd0, dist_reg[8], 6'd0};
		4'd7: n_loc_oh_reg[247] = {8'd0, dist_reg[8], 7'd0};
		4'd8: n_loc_oh_reg[247] = {7'd0, dist_reg[8], 8'd0};
		4'd9: n_loc_oh_reg[247] = {6'd0, dist_reg[8], 9'd0};
		4'd10: n_loc_oh_reg[247] = {5'd0, dist_reg[8], 10'd0};
		4'd11: n_loc_oh_reg[247] = {4'd0, dist_reg[8], 11'd0};
		4'd12: n_loc_oh_reg[247] = {3'd0, dist_reg[8], 12'd0};
		4'd13: n_loc_oh_reg[247] = {2'd0, dist_reg[8], 13'd0};
		4'd14: n_loc_oh_reg[247] = {1'd0, dist_reg[8], 14'd0};
		4'd15: n_loc_oh_reg[247] = {dist_reg[8], 15'd0};
	endcase
	case(loc_reg[248])
		4'd0: n_loc_oh_reg[248] = {15'd0, dist_reg[7]};
		4'd1: n_loc_oh_reg[248] = {14'd0, dist_reg[7], 1'd0};
		4'd2: n_loc_oh_reg[248] = {13'd0, dist_reg[7], 2'd0};
		4'd3: n_loc_oh_reg[248] = {12'd0, dist_reg[7], 3'd0};
		4'd4: n_loc_oh_reg[248] = {11'd0, dist_reg[7], 4'd0};
		4'd5: n_loc_oh_reg[248] = {10'd0, dist_reg[7], 5'd0};
		4'd6: n_loc_oh_reg[248] = {9'd0, dist_reg[7], 6'd0};
		4'd7: n_loc_oh_reg[248] = {8'd0, dist_reg[7], 7'd0};
		4'd8: n_loc_oh_reg[248] = {7'd0, dist_reg[7], 8'd0};
		4'd9: n_loc_oh_reg[248] = {6'd0, dist_reg[7], 9'd0};
		4'd10: n_loc_oh_reg[248] = {5'd0, dist_reg[7], 10'd0};
		4'd11: n_loc_oh_reg[248] = {4'd0, dist_reg[7], 11'd0};
		4'd12: n_loc_oh_reg[248] = {3'd0, dist_reg[7], 12'd0};
		4'd13: n_loc_oh_reg[248] = {2'd0, dist_reg[7], 13'd0};
		4'd14: n_loc_oh_reg[248] = {1'd0, dist_reg[7], 14'd0};
		4'd15: n_loc_oh_reg[248] = {dist_reg[7], 15'd0};
	endcase
	case(loc_reg[249])
		4'd0: n_loc_oh_reg[249] = {15'd0, dist_reg[6]};
		4'd1: n_loc_oh_reg[249] = {14'd0, dist_reg[6], 1'd0};
		4'd2: n_loc_oh_reg[249] = {13'd0, dist_reg[6], 2'd0};
		4'd3: n_loc_oh_reg[249] = {12'd0, dist_reg[6], 3'd0};
		4'd4: n_loc_oh_reg[249] = {11'd0, dist_reg[6], 4'd0};
		4'd5: n_loc_oh_reg[249] = {10'd0, dist_reg[6], 5'd0};
		4'd6: n_loc_oh_reg[249] = {9'd0, dist_reg[6], 6'd0};
		4'd7: n_loc_oh_reg[249] = {8'd0, dist_reg[6], 7'd0};
		4'd8: n_loc_oh_reg[249] = {7'd0, dist_reg[6], 8'd0};
		4'd9: n_loc_oh_reg[249] = {6'd0, dist_reg[6], 9'd0};
		4'd10: n_loc_oh_reg[249] = {5'd0, dist_reg[6], 10'd0};
		4'd11: n_loc_oh_reg[249] = {4'd0, dist_reg[6], 11'd0};
		4'd12: n_loc_oh_reg[249] = {3'd0, dist_reg[6], 12'd0};
		4'd13: n_loc_oh_reg[249] = {2'd0, dist_reg[6], 13'd0};
		4'd14: n_loc_oh_reg[249] = {1'd0, dist_reg[6], 14'd0};
		4'd15: n_loc_oh_reg[249] = {dist_reg[6], 15'd0};
	endcase
	case(loc_reg[250])
		4'd0: n_loc_oh_reg[250] = {15'd0, dist_reg[5]};
		4'd1: n_loc_oh_reg[250] = {14'd0, dist_reg[5], 1'd0};
		4'd2: n_loc_oh_reg[250] = {13'd0, dist_reg[5], 2'd0};
		4'd3: n_loc_oh_reg[250] = {12'd0, dist_reg[5], 3'd0};
		4'd4: n_loc_oh_reg[250] = {11'd0, dist_reg[5], 4'd0};
		4'd5: n_loc_oh_reg[250] = {10'd0, dist_reg[5], 5'd0};
		4'd6: n_loc_oh_reg[250] = {9'd0, dist_reg[5], 6'd0};
		4'd7: n_loc_oh_reg[250] = {8'd0, dist_reg[5], 7'd0};
		4'd8: n_loc_oh_reg[250] = {7'd0, dist_reg[5], 8'd0};
		4'd9: n_loc_oh_reg[250] = {6'd0, dist_reg[5], 9'd0};
		4'd10: n_loc_oh_reg[250] = {5'd0, dist_reg[5], 10'd0};
		4'd11: n_loc_oh_reg[250] = {4'd0, dist_reg[5], 11'd0};
		4'd12: n_loc_oh_reg[250] = {3'd0, dist_reg[5], 12'd0};
		4'd13: n_loc_oh_reg[250] = {2'd0, dist_reg[5], 13'd0};
		4'd14: n_loc_oh_reg[250] = {1'd0, dist_reg[5], 14'd0};
		4'd15: n_loc_oh_reg[250] = {dist_reg[5], 15'd0};
	endcase
	case(loc_reg[251])
		4'd0: n_loc_oh_reg[251] = {15'd0, dist_reg[4]};
		4'd1: n_loc_oh_reg[251] = {14'd0, dist_reg[4], 1'd0};
		4'd2: n_loc_oh_reg[251] = {13'd0, dist_reg[4], 2'd0};
		4'd3: n_loc_oh_reg[251] = {12'd0, dist_reg[4], 3'd0};
		4'd4: n_loc_oh_reg[251] = {11'd0, dist_reg[4], 4'd0};
		4'd5: n_loc_oh_reg[251] = {10'd0, dist_reg[4], 5'd0};
		4'd6: n_loc_oh_reg[251] = {9'd0, dist_reg[4], 6'd0};
		4'd7: n_loc_oh_reg[251] = {8'd0, dist_reg[4], 7'd0};
		4'd8: n_loc_oh_reg[251] = {7'd0, dist_reg[4], 8'd0};
		4'd9: n_loc_oh_reg[251] = {6'd0, dist_reg[4], 9'd0};
		4'd10: n_loc_oh_reg[251] = {5'd0, dist_reg[4], 10'd0};
		4'd11: n_loc_oh_reg[251] = {4'd0, dist_reg[4], 11'd0};
		4'd12: n_loc_oh_reg[251] = {3'd0, dist_reg[4], 12'd0};
		4'd13: n_loc_oh_reg[251] = {2'd0, dist_reg[4], 13'd0};
		4'd14: n_loc_oh_reg[251] = {1'd0, dist_reg[4], 14'd0};
		4'd15: n_loc_oh_reg[251] = {dist_reg[4], 15'd0};
	endcase
	case(loc_reg[252])
		4'd0: n_loc_oh_reg[252] = {15'd0, dist_reg[3]};
		4'd1: n_loc_oh_reg[252] = {14'd0, dist_reg[3], 1'd0};
		4'd2: n_loc_oh_reg[252] = {13'd0, dist_reg[3], 2'd0};
		4'd3: n_loc_oh_reg[252] = {12'd0, dist_reg[3], 3'd0};
		4'd4: n_loc_oh_reg[252] = {11'd0, dist_reg[3], 4'd0};
		4'd5: n_loc_oh_reg[252] = {10'd0, dist_reg[3], 5'd0};
		4'd6: n_loc_oh_reg[252] = {9'd0, dist_reg[3], 6'd0};
		4'd7: n_loc_oh_reg[252] = {8'd0, dist_reg[3], 7'd0};
		4'd8: n_loc_oh_reg[252] = {7'd0, dist_reg[3], 8'd0};
		4'd9: n_loc_oh_reg[252] = {6'd0, dist_reg[3], 9'd0};
		4'd10: n_loc_oh_reg[252] = {5'd0, dist_reg[3], 10'd0};
		4'd11: n_loc_oh_reg[252] = {4'd0, dist_reg[3], 11'd0};
		4'd12: n_loc_oh_reg[252] = {3'd0, dist_reg[3], 12'd0};
		4'd13: n_loc_oh_reg[252] = {2'd0, dist_reg[3], 13'd0};
		4'd14: n_loc_oh_reg[252] = {1'd0, dist_reg[3], 14'd0};
		4'd15: n_loc_oh_reg[252] = {dist_reg[3], 15'd0};
	endcase
	case(loc_reg[253])
		4'd0: n_loc_oh_reg[253] = {15'd0, dist_reg[2]};
		4'd1: n_loc_oh_reg[253] = {14'd0, dist_reg[2], 1'd0};
		4'd2: n_loc_oh_reg[253] = {13'd0, dist_reg[2], 2'd0};
		4'd3: n_loc_oh_reg[253] = {12'd0, dist_reg[2], 3'd0};
		4'd4: n_loc_oh_reg[253] = {11'd0, dist_reg[2], 4'd0};
		4'd5: n_loc_oh_reg[253] = {10'd0, dist_reg[2], 5'd0};
		4'd6: n_loc_oh_reg[253] = {9'd0, dist_reg[2], 6'd0};
		4'd7: n_loc_oh_reg[253] = {8'd0, dist_reg[2], 7'd0};
		4'd8: n_loc_oh_reg[253] = {7'd0, dist_reg[2], 8'd0};
		4'd9: n_loc_oh_reg[253] = {6'd0, dist_reg[2], 9'd0};
		4'd10: n_loc_oh_reg[253] = {5'd0, dist_reg[2], 10'd0};
		4'd11: n_loc_oh_reg[253] = {4'd0, dist_reg[2], 11'd0};
		4'd12: n_loc_oh_reg[253] = {3'd0, dist_reg[2], 12'd0};
		4'd13: n_loc_oh_reg[253] = {2'd0, dist_reg[2], 13'd0};
		4'd14: n_loc_oh_reg[253] = {1'd0, dist_reg[2], 14'd0};
		4'd15: n_loc_oh_reg[253] = {dist_reg[2], 15'd0};
	endcase
	case(loc_reg[254])
		4'd0: n_loc_oh_reg[254] = {15'd0, dist_reg[1]};
		4'd1: n_loc_oh_reg[254] = {14'd0, dist_reg[1], 1'd0};
		4'd2: n_loc_oh_reg[254] = {13'd0, dist_reg[1], 2'd0};
		4'd3: n_loc_oh_reg[254] = {12'd0, dist_reg[1], 3'd0};
		4'd4: n_loc_oh_reg[254] = {11'd0, dist_reg[1], 4'd0};
		4'd5: n_loc_oh_reg[254] = {10'd0, dist_reg[1], 5'd0};
		4'd6: n_loc_oh_reg[254] = {9'd0, dist_reg[1], 6'd0};
		4'd7: n_loc_oh_reg[254] = {8'd0, dist_reg[1], 7'd0};
		4'd8: n_loc_oh_reg[254] = {7'd0, dist_reg[1], 8'd0};
		4'd9: n_loc_oh_reg[254] = {6'd0, dist_reg[1], 9'd0};
		4'd10: n_loc_oh_reg[254] = {5'd0, dist_reg[1], 10'd0};
		4'd11: n_loc_oh_reg[254] = {4'd0, dist_reg[1], 11'd0};
		4'd12: n_loc_oh_reg[254] = {3'd0, dist_reg[1], 12'd0};
		4'd13: n_loc_oh_reg[254] = {2'd0, dist_reg[1], 13'd0};
		4'd14: n_loc_oh_reg[254] = {1'd0, dist_reg[1], 14'd0};
		4'd15: n_loc_oh_reg[254] = {dist_reg[1], 15'd0};
	endcase
	case(loc_reg[255])
		4'd0: n_loc_oh_reg[255] = {15'd0, dist_reg[0]};
		4'd1: n_loc_oh_reg[255] = {14'd0, dist_reg[0], 1'd0};
		4'd2: n_loc_oh_reg[255] = {13'd0, dist_reg[0], 2'd0};
		4'd3: n_loc_oh_reg[255] = {12'd0, dist_reg[0], 3'd0};
		4'd4: n_loc_oh_reg[255] = {11'd0, dist_reg[0], 4'd0};
		4'd5: n_loc_oh_reg[255] = {10'd0, dist_reg[0], 5'd0};
		4'd6: n_loc_oh_reg[255] = {9'd0, dist_reg[0], 6'd0};
		4'd7: n_loc_oh_reg[255] = {8'd0, dist_reg[0], 7'd0};
		4'd8: n_loc_oh_reg[255] = {7'd0, dist_reg[0], 8'd0};
		4'd9: n_loc_oh_reg[255] = {6'd0, dist_reg[0], 9'd0};
		4'd10: n_loc_oh_reg[255] = {5'd0, dist_reg[0], 10'd0};
		4'd11: n_loc_oh_reg[255] = {4'd0, dist_reg[0], 11'd0};
		4'd12: n_loc_oh_reg[255] = {3'd0, dist_reg[0], 12'd0};
		4'd13: n_loc_oh_reg[255] = {2'd0, dist_reg[0], 13'd0};
		4'd14: n_loc_oh_reg[255] = {1'd0, dist_reg[0], 14'd0};
		4'd15: n_loc_oh_reg[255] = {dist_reg[0], 15'd0};
	endcase
end

// COMB2: get dsum_reg
always@* begin
    n_dsum_reg[0] = loc_oh_reg[0][0] + loc_oh_reg[1][0] + loc_oh_reg[2][0] + loc_oh_reg[3][0] + loc_oh_reg[4][0] + loc_oh_reg[5][0] + loc_oh_reg[6][0] + loc_oh_reg[7][0] + loc_oh_reg[8][0] + loc_oh_reg[9][0] + loc_oh_reg[10][0] + loc_oh_reg[11][0] + loc_oh_reg[12][0] + loc_oh_reg[13][0] + loc_oh_reg[14][0] + loc_oh_reg[15][0] + loc_oh_reg[16][0] + loc_oh_reg[17][0] + loc_oh_reg[18][0] + loc_oh_reg[19][0] + loc_oh_reg[20][0] + loc_oh_reg[21][0] + loc_oh_reg[22][0] + loc_oh_reg[23][0] + loc_oh_reg[24][0] + loc_oh_reg[25][0] + loc_oh_reg[26][0] + loc_oh_reg[27][0] + loc_oh_reg[28][0] + loc_oh_reg[29][0] + loc_oh_reg[30][0] + loc_oh_reg[31][0];
    n_dsum_reg[1] = loc_oh_reg[32][0] + loc_oh_reg[33][0] + loc_oh_reg[34][0] + loc_oh_reg[35][0] + loc_oh_reg[36][0] + loc_oh_reg[37][0] + loc_oh_reg[38][0] + loc_oh_reg[39][0] + loc_oh_reg[40][0] + loc_oh_reg[41][0] + loc_oh_reg[42][0] + loc_oh_reg[43][0] + loc_oh_reg[44][0] + loc_oh_reg[45][0] + loc_oh_reg[46][0] + loc_oh_reg[47][0] + loc_oh_reg[48][0] + loc_oh_reg[49][0] + loc_oh_reg[50][0] + loc_oh_reg[51][0] + loc_oh_reg[52][0] + loc_oh_reg[53][0] + loc_oh_reg[54][0] + loc_oh_reg[55][0] + loc_oh_reg[56][0] + loc_oh_reg[57][0] + loc_oh_reg[58][0] + loc_oh_reg[59][0] + loc_oh_reg[60][0] + loc_oh_reg[61][0] + loc_oh_reg[62][0] + loc_oh_reg[63][0];
    n_dsum_reg[2] = loc_oh_reg[64][0] + loc_oh_reg[65][0] + loc_oh_reg[66][0] + loc_oh_reg[67][0] + loc_oh_reg[68][0] + loc_oh_reg[69][0] + loc_oh_reg[70][0] + loc_oh_reg[71][0] + loc_oh_reg[72][0] + loc_oh_reg[73][0] + loc_oh_reg[74][0] + loc_oh_reg[75][0] + loc_oh_reg[76][0] + loc_oh_reg[77][0] + loc_oh_reg[78][0] + loc_oh_reg[79][0] + loc_oh_reg[80][0] + loc_oh_reg[81][0] + loc_oh_reg[82][0] + loc_oh_reg[83][0] + loc_oh_reg[84][0] + loc_oh_reg[85][0] + loc_oh_reg[86][0] + loc_oh_reg[87][0] + loc_oh_reg[88][0] + loc_oh_reg[89][0] + loc_oh_reg[90][0] + loc_oh_reg[91][0] + loc_oh_reg[92][0] + loc_oh_reg[93][0] + loc_oh_reg[94][0] + loc_oh_reg[95][0];
    n_dsum_reg[3] = loc_oh_reg[96][0] + loc_oh_reg[97][0] + loc_oh_reg[98][0] + loc_oh_reg[99][0] + loc_oh_reg[100][0] + loc_oh_reg[101][0] + loc_oh_reg[102][0] + loc_oh_reg[103][0] + loc_oh_reg[104][0] + loc_oh_reg[105][0] + loc_oh_reg[106][0] + loc_oh_reg[107][0] + loc_oh_reg[108][0] + loc_oh_reg[109][0] + loc_oh_reg[110][0] + loc_oh_reg[111][0] + loc_oh_reg[112][0] + loc_oh_reg[113][0] + loc_oh_reg[114][0] + loc_oh_reg[115][0] + loc_oh_reg[116][0] + loc_oh_reg[117][0] + loc_oh_reg[118][0] + loc_oh_reg[119][0] + loc_oh_reg[120][0] + loc_oh_reg[121][0] + loc_oh_reg[122][0] + loc_oh_reg[123][0] + loc_oh_reg[124][0] + loc_oh_reg[125][0] + loc_oh_reg[126][0] + loc_oh_reg[127][0];
    n_dsum_reg[4] = loc_oh_reg[128][0] + loc_oh_reg[129][0] + loc_oh_reg[130][0] + loc_oh_reg[131][0] + loc_oh_reg[132][0] + loc_oh_reg[133][0] + loc_oh_reg[134][0] + loc_oh_reg[135][0] + loc_oh_reg[136][0] + loc_oh_reg[137][0] + loc_oh_reg[138][0] + loc_oh_reg[139][0] + loc_oh_reg[140][0] + loc_oh_reg[141][0] + loc_oh_reg[142][0] + loc_oh_reg[143][0] + loc_oh_reg[144][0] + loc_oh_reg[145][0] + loc_oh_reg[146][0] + loc_oh_reg[147][0] + loc_oh_reg[148][0] + loc_oh_reg[149][0] + loc_oh_reg[150][0] + loc_oh_reg[151][0] + loc_oh_reg[152][0] + loc_oh_reg[153][0] + loc_oh_reg[154][0] + loc_oh_reg[155][0] + loc_oh_reg[156][0] + loc_oh_reg[157][0] + loc_oh_reg[158][0] + loc_oh_reg[159][0];
    n_dsum_reg[5] = loc_oh_reg[160][0] + loc_oh_reg[161][0] + loc_oh_reg[162][0] + loc_oh_reg[163][0] + loc_oh_reg[164][0] + loc_oh_reg[165][0] + loc_oh_reg[166][0] + loc_oh_reg[167][0] + loc_oh_reg[168][0] + loc_oh_reg[169][0] + loc_oh_reg[170][0] + loc_oh_reg[171][0] + loc_oh_reg[172][0] + loc_oh_reg[173][0] + loc_oh_reg[174][0] + loc_oh_reg[175][0] + loc_oh_reg[176][0] + loc_oh_reg[177][0] + loc_oh_reg[178][0] + loc_oh_reg[179][0] + loc_oh_reg[180][0] + loc_oh_reg[181][0] + loc_oh_reg[182][0] + loc_oh_reg[183][0] + loc_oh_reg[184][0] + loc_oh_reg[185][0] + loc_oh_reg[186][0] + loc_oh_reg[187][0] + loc_oh_reg[188][0] + loc_oh_reg[189][0] + loc_oh_reg[190][0] + loc_oh_reg[191][0];
    n_dsum_reg[6] = loc_oh_reg[192][0] + loc_oh_reg[193][0] + loc_oh_reg[194][0] + loc_oh_reg[195][0] + loc_oh_reg[196][0] + loc_oh_reg[197][0] + loc_oh_reg[198][0] + loc_oh_reg[199][0] + loc_oh_reg[200][0] + loc_oh_reg[201][0] + loc_oh_reg[202][0] + loc_oh_reg[203][0] + loc_oh_reg[204][0] + loc_oh_reg[205][0] + loc_oh_reg[206][0] + loc_oh_reg[207][0] + loc_oh_reg[208][0] + loc_oh_reg[209][0] + loc_oh_reg[210][0] + loc_oh_reg[211][0] + loc_oh_reg[212][0] + loc_oh_reg[213][0] + loc_oh_reg[214][0] + loc_oh_reg[215][0] + loc_oh_reg[216][0] + loc_oh_reg[217][0] + loc_oh_reg[218][0] + loc_oh_reg[219][0] + loc_oh_reg[220][0] + loc_oh_reg[221][0] + loc_oh_reg[222][0] + loc_oh_reg[223][0];
    n_dsum_reg[7] = loc_oh_reg[224][0] + loc_oh_reg[225][0] + loc_oh_reg[226][0] + loc_oh_reg[227][0] + loc_oh_reg[228][0] + loc_oh_reg[229][0] + loc_oh_reg[230][0] + loc_oh_reg[231][0] + loc_oh_reg[232][0] + loc_oh_reg[233][0] + loc_oh_reg[234][0] + loc_oh_reg[235][0] + loc_oh_reg[236][0] + loc_oh_reg[237][0] + loc_oh_reg[238][0] + loc_oh_reg[239][0] + loc_oh_reg[240][0] + loc_oh_reg[241][0] + loc_oh_reg[242][0] + loc_oh_reg[243][0] + loc_oh_reg[244][0] + loc_oh_reg[245][0] + loc_oh_reg[246][0] + loc_oh_reg[247][0] + loc_oh_reg[248][0] + loc_oh_reg[249][0] + loc_oh_reg[250][0] + loc_oh_reg[251][0] + loc_oh_reg[252][0] + loc_oh_reg[253][0] + loc_oh_reg[254][0] + loc_oh_reg[255][0];

    n_dsum_reg[8] = loc_oh_reg[0][1] + loc_oh_reg[1][1] + loc_oh_reg[2][1] + loc_oh_reg[3][1] + loc_oh_reg[4][1] + loc_oh_reg[5][1] + loc_oh_reg[6][1] + loc_oh_reg[7][1] + loc_oh_reg[8][1] + loc_oh_reg[9][1] + loc_oh_reg[10][1] + loc_oh_reg[11][1] + loc_oh_reg[12][1] + loc_oh_reg[13][1] + loc_oh_reg[14][1] + loc_oh_reg[15][1] + loc_oh_reg[16][1] + loc_oh_reg[17][1] + loc_oh_reg[18][1] + loc_oh_reg[19][1] + loc_oh_reg[20][1] + loc_oh_reg[21][1] + loc_oh_reg[22][1] + loc_oh_reg[23][1] + loc_oh_reg[24][1] + loc_oh_reg[25][1] + loc_oh_reg[26][1] + loc_oh_reg[27][1] + loc_oh_reg[28][1] + loc_oh_reg[29][1] + loc_oh_reg[30][1] + loc_oh_reg[31][1];
    n_dsum_reg[9] = loc_oh_reg[32][1] + loc_oh_reg[33][1] + loc_oh_reg[34][1] + loc_oh_reg[35][1] + loc_oh_reg[36][1] + loc_oh_reg[37][1] + loc_oh_reg[38][1] + loc_oh_reg[39][1] + loc_oh_reg[40][1] + loc_oh_reg[41][1] + loc_oh_reg[42][1] + loc_oh_reg[43][1] + loc_oh_reg[44][1] + loc_oh_reg[45][1] + loc_oh_reg[46][1] + loc_oh_reg[47][1] + loc_oh_reg[48][1] + loc_oh_reg[49][1] + loc_oh_reg[50][1] + loc_oh_reg[51][1] + loc_oh_reg[52][1] + loc_oh_reg[53][1] + loc_oh_reg[54][1] + loc_oh_reg[55][1] + loc_oh_reg[56][1] + loc_oh_reg[57][1] + loc_oh_reg[58][1] + loc_oh_reg[59][1] + loc_oh_reg[60][1] + loc_oh_reg[61][1] + loc_oh_reg[62][1] + loc_oh_reg[63][1];
    n_dsum_reg[10] = loc_oh_reg[64][1] + loc_oh_reg[65][1] + loc_oh_reg[66][1] + loc_oh_reg[67][1] + loc_oh_reg[68][1] + loc_oh_reg[69][1] + loc_oh_reg[70][1] + loc_oh_reg[71][1] + loc_oh_reg[72][1] + loc_oh_reg[73][1] + loc_oh_reg[74][1] + loc_oh_reg[75][1] + loc_oh_reg[76][1] + loc_oh_reg[77][1] + loc_oh_reg[78][1] + loc_oh_reg[79][1] + loc_oh_reg[80][1] + loc_oh_reg[81][1] + loc_oh_reg[82][1] + loc_oh_reg[83][1] + loc_oh_reg[84][1] + loc_oh_reg[85][1] + loc_oh_reg[86][1] + loc_oh_reg[87][1] + loc_oh_reg[88][1] + loc_oh_reg[89][1] + loc_oh_reg[90][1] + loc_oh_reg[91][1] + loc_oh_reg[92][1] + loc_oh_reg[93][1] + loc_oh_reg[94][1] + loc_oh_reg[95][1];
    n_dsum_reg[11] = loc_oh_reg[96][1] + loc_oh_reg[97][1] + loc_oh_reg[98][1] + loc_oh_reg[99][1] + loc_oh_reg[100][1] + loc_oh_reg[101][1] + loc_oh_reg[102][1] + loc_oh_reg[103][1] + loc_oh_reg[104][1] + loc_oh_reg[105][1] + loc_oh_reg[106][1] + loc_oh_reg[107][1] + loc_oh_reg[108][1] + loc_oh_reg[109][1] + loc_oh_reg[110][1] + loc_oh_reg[111][1] + loc_oh_reg[112][1] + loc_oh_reg[113][1] + loc_oh_reg[114][1] + loc_oh_reg[115][1] + loc_oh_reg[116][1] + loc_oh_reg[117][1] + loc_oh_reg[118][1] + loc_oh_reg[119][1] + loc_oh_reg[120][1] + loc_oh_reg[121][1] + loc_oh_reg[122][1] + loc_oh_reg[123][1] + loc_oh_reg[124][1] + loc_oh_reg[125][1] + loc_oh_reg[126][1] + loc_oh_reg[127][1];
    n_dsum_reg[12] = loc_oh_reg[128][1] + loc_oh_reg[129][1] + loc_oh_reg[130][1] + loc_oh_reg[131][1] + loc_oh_reg[132][1] + loc_oh_reg[133][1] + loc_oh_reg[134][1] + loc_oh_reg[135][1] + loc_oh_reg[136][1] + loc_oh_reg[137][1] + loc_oh_reg[138][1] + loc_oh_reg[139][1] + loc_oh_reg[140][1] + loc_oh_reg[141][1] + loc_oh_reg[142][1] + loc_oh_reg[143][1] + loc_oh_reg[144][1] + loc_oh_reg[145][1] + loc_oh_reg[146][1] + loc_oh_reg[147][1] + loc_oh_reg[148][1] + loc_oh_reg[149][1] + loc_oh_reg[150][1] + loc_oh_reg[151][1] + loc_oh_reg[152][1] + loc_oh_reg[153][1] + loc_oh_reg[154][1] + loc_oh_reg[155][1] + loc_oh_reg[156][1] + loc_oh_reg[157][1] + loc_oh_reg[158][1] + loc_oh_reg[159][1];
    n_dsum_reg[13] = loc_oh_reg[160][1] + loc_oh_reg[161][1] + loc_oh_reg[162][1] + loc_oh_reg[163][1] + loc_oh_reg[164][1] + loc_oh_reg[165][1] + loc_oh_reg[166][1] + loc_oh_reg[167][1] + loc_oh_reg[168][1] + loc_oh_reg[169][1] + loc_oh_reg[170][1] + loc_oh_reg[171][1] + loc_oh_reg[172][1] + loc_oh_reg[173][1] + loc_oh_reg[174][1] + loc_oh_reg[175][1] + loc_oh_reg[176][1] + loc_oh_reg[177][1] + loc_oh_reg[178][1] + loc_oh_reg[179][1] + loc_oh_reg[180][1] + loc_oh_reg[181][1] + loc_oh_reg[182][1] + loc_oh_reg[183][1] + loc_oh_reg[184][1] + loc_oh_reg[185][1] + loc_oh_reg[186][1] + loc_oh_reg[187][1] + loc_oh_reg[188][1] + loc_oh_reg[189][1] + loc_oh_reg[190][1] + loc_oh_reg[191][1];
    n_dsum_reg[14] = loc_oh_reg[192][1] + loc_oh_reg[193][1] + loc_oh_reg[194][1] + loc_oh_reg[195][1] + loc_oh_reg[196][1] + loc_oh_reg[197][1] + loc_oh_reg[198][1] + loc_oh_reg[199][1] + loc_oh_reg[200][1] + loc_oh_reg[201][1] + loc_oh_reg[202][1] + loc_oh_reg[203][1] + loc_oh_reg[204][1] + loc_oh_reg[205][1] + loc_oh_reg[206][1] + loc_oh_reg[207][1] + loc_oh_reg[208][1] + loc_oh_reg[209][1] + loc_oh_reg[210][1] + loc_oh_reg[211][1] + loc_oh_reg[212][1] + loc_oh_reg[213][1] + loc_oh_reg[214][1] + loc_oh_reg[215][1] + loc_oh_reg[216][1] + loc_oh_reg[217][1] + loc_oh_reg[218][1] + loc_oh_reg[219][1] + loc_oh_reg[220][1] + loc_oh_reg[221][1] + loc_oh_reg[222][1] + loc_oh_reg[223][1];
    n_dsum_reg[15] = loc_oh_reg[224][1] + loc_oh_reg[225][1] + loc_oh_reg[226][1] + loc_oh_reg[227][1] + loc_oh_reg[228][1] + loc_oh_reg[229][1] + loc_oh_reg[230][1] + loc_oh_reg[231][1] + loc_oh_reg[232][1] + loc_oh_reg[233][1] + loc_oh_reg[234][1] + loc_oh_reg[235][1] + loc_oh_reg[236][1] + loc_oh_reg[237][1] + loc_oh_reg[238][1] + loc_oh_reg[239][1] + loc_oh_reg[240][1] + loc_oh_reg[241][1] + loc_oh_reg[242][1] + loc_oh_reg[243][1] + loc_oh_reg[244][1] + loc_oh_reg[245][1] + loc_oh_reg[246][1] + loc_oh_reg[247][1] + loc_oh_reg[248][1] + loc_oh_reg[249][1] + loc_oh_reg[250][1] + loc_oh_reg[251][1] + loc_oh_reg[252][1] + loc_oh_reg[253][1] + loc_oh_reg[254][1] + loc_oh_reg[255][1];

    n_dsum_reg[16] = loc_oh_reg[0][2] + loc_oh_reg[1][2] + loc_oh_reg[2][2] + loc_oh_reg[3][2] + loc_oh_reg[4][2] + loc_oh_reg[5][2] + loc_oh_reg[6][2] + loc_oh_reg[7][2] + loc_oh_reg[8][2] + loc_oh_reg[9][2] + loc_oh_reg[10][2] + loc_oh_reg[11][2] + loc_oh_reg[12][2] + loc_oh_reg[13][2] + loc_oh_reg[14][2] + loc_oh_reg[15][2] + loc_oh_reg[16][2] + loc_oh_reg[17][2] + loc_oh_reg[18][2] + loc_oh_reg[19][2] + loc_oh_reg[20][2] + loc_oh_reg[21][2] + loc_oh_reg[22][2] + loc_oh_reg[23][2] + loc_oh_reg[24][2] + loc_oh_reg[25][2] + loc_oh_reg[26][2] + loc_oh_reg[27][2] + loc_oh_reg[28][2] + loc_oh_reg[29][2] + loc_oh_reg[30][2] + loc_oh_reg[31][2];
    n_dsum_reg[17] = loc_oh_reg[32][2] + loc_oh_reg[33][2] + loc_oh_reg[34][2] + loc_oh_reg[35][2] + loc_oh_reg[36][2] + loc_oh_reg[37][2] + loc_oh_reg[38][2] + loc_oh_reg[39][2] + loc_oh_reg[40][2] + loc_oh_reg[41][2] + loc_oh_reg[42][2] + loc_oh_reg[43][2] + loc_oh_reg[44][2] + loc_oh_reg[45][2] + loc_oh_reg[46][2] + loc_oh_reg[47][2] + loc_oh_reg[48][2] + loc_oh_reg[49][2] + loc_oh_reg[50][2] + loc_oh_reg[51][2] + loc_oh_reg[52][2] + loc_oh_reg[53][2] + loc_oh_reg[54][2] + loc_oh_reg[55][2] + loc_oh_reg[56][2] + loc_oh_reg[57][2] + loc_oh_reg[58][2] + loc_oh_reg[59][2] + loc_oh_reg[60][2] + loc_oh_reg[61][2] + loc_oh_reg[62][2] + loc_oh_reg[63][2];
    n_dsum_reg[18] = loc_oh_reg[64][2] + loc_oh_reg[65][2] + loc_oh_reg[66][2] + loc_oh_reg[67][2] + loc_oh_reg[68][2] + loc_oh_reg[69][2] + loc_oh_reg[70][2] + loc_oh_reg[71][2] + loc_oh_reg[72][2] + loc_oh_reg[73][2] + loc_oh_reg[74][2] + loc_oh_reg[75][2] + loc_oh_reg[76][2] + loc_oh_reg[77][2] + loc_oh_reg[78][2] + loc_oh_reg[79][2] + loc_oh_reg[80][2] + loc_oh_reg[81][2] + loc_oh_reg[82][2] + loc_oh_reg[83][2] + loc_oh_reg[84][2] + loc_oh_reg[85][2] + loc_oh_reg[86][2] + loc_oh_reg[87][2] + loc_oh_reg[88][2] + loc_oh_reg[89][2] + loc_oh_reg[90][2] + loc_oh_reg[91][2] + loc_oh_reg[92][2] + loc_oh_reg[93][2] + loc_oh_reg[94][2] + loc_oh_reg[95][2];
    n_dsum_reg[19] = loc_oh_reg[96][2] + loc_oh_reg[97][2] + loc_oh_reg[98][2] + loc_oh_reg[99][2] + loc_oh_reg[100][2] + loc_oh_reg[101][2] + loc_oh_reg[102][2] + loc_oh_reg[103][2] + loc_oh_reg[104][2] + loc_oh_reg[105][2] + loc_oh_reg[106][2] + loc_oh_reg[107][2] + loc_oh_reg[108][2] + loc_oh_reg[109][2] + loc_oh_reg[110][2] + loc_oh_reg[111][2] + loc_oh_reg[112][2] + loc_oh_reg[113][2] + loc_oh_reg[114][2] + loc_oh_reg[115][2] + loc_oh_reg[116][2] + loc_oh_reg[117][2] + loc_oh_reg[118][2] + loc_oh_reg[119][2] + loc_oh_reg[120][2] + loc_oh_reg[121][2] + loc_oh_reg[122][2] + loc_oh_reg[123][2] + loc_oh_reg[124][2] + loc_oh_reg[125][2] + loc_oh_reg[126][2] + loc_oh_reg[127][2];
    n_dsum_reg[20] = loc_oh_reg[128][2] + loc_oh_reg[129][2] + loc_oh_reg[130][2] + loc_oh_reg[131][2] + loc_oh_reg[132][2] + loc_oh_reg[133][2] + loc_oh_reg[134][2] + loc_oh_reg[135][2] + loc_oh_reg[136][2] + loc_oh_reg[137][2] + loc_oh_reg[138][2] + loc_oh_reg[139][2] + loc_oh_reg[140][2] + loc_oh_reg[141][2] + loc_oh_reg[142][2] + loc_oh_reg[143][2] + loc_oh_reg[144][2] + loc_oh_reg[145][2] + loc_oh_reg[146][2] + loc_oh_reg[147][2] + loc_oh_reg[148][2] + loc_oh_reg[149][2] + loc_oh_reg[150][2] + loc_oh_reg[151][2] + loc_oh_reg[152][2] + loc_oh_reg[153][2] + loc_oh_reg[154][2] + loc_oh_reg[155][2] + loc_oh_reg[156][2] + loc_oh_reg[157][2] + loc_oh_reg[158][2] + loc_oh_reg[159][2];
    n_dsum_reg[21] = loc_oh_reg[160][2] + loc_oh_reg[161][2] + loc_oh_reg[162][2] + loc_oh_reg[163][2] + loc_oh_reg[164][2] + loc_oh_reg[165][2] + loc_oh_reg[166][2] + loc_oh_reg[167][2] + loc_oh_reg[168][2] + loc_oh_reg[169][2] + loc_oh_reg[170][2] + loc_oh_reg[171][2] + loc_oh_reg[172][2] + loc_oh_reg[173][2] + loc_oh_reg[174][2] + loc_oh_reg[175][2] + loc_oh_reg[176][2] + loc_oh_reg[177][2] + loc_oh_reg[178][2] + loc_oh_reg[179][2] + loc_oh_reg[180][2] + loc_oh_reg[181][2] + loc_oh_reg[182][2] + loc_oh_reg[183][2] + loc_oh_reg[184][2] + loc_oh_reg[185][2] + loc_oh_reg[186][2] + loc_oh_reg[187][2] + loc_oh_reg[188][2] + loc_oh_reg[189][2] + loc_oh_reg[190][2] + loc_oh_reg[191][2];
    n_dsum_reg[22] = loc_oh_reg[192][2] + loc_oh_reg[193][2] + loc_oh_reg[194][2] + loc_oh_reg[195][2] + loc_oh_reg[196][2] + loc_oh_reg[197][2] + loc_oh_reg[198][2] + loc_oh_reg[199][2] + loc_oh_reg[200][2] + loc_oh_reg[201][2] + loc_oh_reg[202][2] + loc_oh_reg[203][2] + loc_oh_reg[204][2] + loc_oh_reg[205][2] + loc_oh_reg[206][2] + loc_oh_reg[207][2] + loc_oh_reg[208][2] + loc_oh_reg[209][2] + loc_oh_reg[210][2] + loc_oh_reg[211][2] + loc_oh_reg[212][2] + loc_oh_reg[213][2] + loc_oh_reg[214][2] + loc_oh_reg[215][2] + loc_oh_reg[216][2] + loc_oh_reg[217][2] + loc_oh_reg[218][2] + loc_oh_reg[219][2] + loc_oh_reg[220][2] + loc_oh_reg[221][2] + loc_oh_reg[222][2] + loc_oh_reg[223][2];
    n_dsum_reg[23] = loc_oh_reg[224][2] + loc_oh_reg[225][2] + loc_oh_reg[226][2] + loc_oh_reg[227][2] + loc_oh_reg[228][2] + loc_oh_reg[229][2] + loc_oh_reg[230][2] + loc_oh_reg[231][2] + loc_oh_reg[232][2] + loc_oh_reg[233][2] + loc_oh_reg[234][2] + loc_oh_reg[235][2] + loc_oh_reg[236][2] + loc_oh_reg[237][2] + loc_oh_reg[238][2] + loc_oh_reg[239][2] + loc_oh_reg[240][2] + loc_oh_reg[241][2] + loc_oh_reg[242][2] + loc_oh_reg[243][2] + loc_oh_reg[244][2] + loc_oh_reg[245][2] + loc_oh_reg[246][2] + loc_oh_reg[247][2] + loc_oh_reg[248][2] + loc_oh_reg[249][2] + loc_oh_reg[250][2] + loc_oh_reg[251][2] + loc_oh_reg[252][2] + loc_oh_reg[253][2] + loc_oh_reg[254][2] + loc_oh_reg[255][2];

    n_dsum_reg[24] = loc_oh_reg[0][3] + loc_oh_reg[1][3] + loc_oh_reg[2][3] + loc_oh_reg[3][3] + loc_oh_reg[4][3] + loc_oh_reg[5][3] + loc_oh_reg[6][3] + loc_oh_reg[7][3] + loc_oh_reg[8][3] + loc_oh_reg[9][3] + loc_oh_reg[10][3] + loc_oh_reg[11][3] + loc_oh_reg[12][3] + loc_oh_reg[13][3] + loc_oh_reg[14][3] + loc_oh_reg[15][3] + loc_oh_reg[16][3] + loc_oh_reg[17][3] + loc_oh_reg[18][3] + loc_oh_reg[19][3] + loc_oh_reg[20][3] + loc_oh_reg[21][3] + loc_oh_reg[22][3] + loc_oh_reg[23][3] + loc_oh_reg[24][3] + loc_oh_reg[25][3] + loc_oh_reg[26][3] + loc_oh_reg[27][3] + loc_oh_reg[28][3] + loc_oh_reg[29][3] + loc_oh_reg[30][3] + loc_oh_reg[31][3];
    n_dsum_reg[25] = loc_oh_reg[32][3] + loc_oh_reg[33][3] + loc_oh_reg[34][3] + loc_oh_reg[35][3] + loc_oh_reg[36][3] + loc_oh_reg[37][3] + loc_oh_reg[38][3] + loc_oh_reg[39][3] + loc_oh_reg[40][3] + loc_oh_reg[41][3] + loc_oh_reg[42][3] + loc_oh_reg[43][3] + loc_oh_reg[44][3] + loc_oh_reg[45][3] + loc_oh_reg[46][3] + loc_oh_reg[47][3] + loc_oh_reg[48][3] + loc_oh_reg[49][3] + loc_oh_reg[50][3] + loc_oh_reg[51][3] + loc_oh_reg[52][3] + loc_oh_reg[53][3] + loc_oh_reg[54][3] + loc_oh_reg[55][3] + loc_oh_reg[56][3] + loc_oh_reg[57][3] + loc_oh_reg[58][3] + loc_oh_reg[59][3] + loc_oh_reg[60][3] + loc_oh_reg[61][3] + loc_oh_reg[62][3] + loc_oh_reg[63][3];
    n_dsum_reg[26] = loc_oh_reg[64][3] + loc_oh_reg[65][3] + loc_oh_reg[66][3] + loc_oh_reg[67][3] + loc_oh_reg[68][3] + loc_oh_reg[69][3] + loc_oh_reg[70][3] + loc_oh_reg[71][3] + loc_oh_reg[72][3] + loc_oh_reg[73][3] + loc_oh_reg[74][3] + loc_oh_reg[75][3] + loc_oh_reg[76][3] + loc_oh_reg[77][3] + loc_oh_reg[78][3] + loc_oh_reg[79][3] + loc_oh_reg[80][3] + loc_oh_reg[81][3] + loc_oh_reg[82][3] + loc_oh_reg[83][3] + loc_oh_reg[84][3] + loc_oh_reg[85][3] + loc_oh_reg[86][3] + loc_oh_reg[87][3] + loc_oh_reg[88][3] + loc_oh_reg[89][3] + loc_oh_reg[90][3] + loc_oh_reg[91][3] + loc_oh_reg[92][3] + loc_oh_reg[93][3] + loc_oh_reg[94][3] + loc_oh_reg[95][3];
    n_dsum_reg[27] = loc_oh_reg[96][3] + loc_oh_reg[97][3] + loc_oh_reg[98][3] + loc_oh_reg[99][3] + loc_oh_reg[100][3] + loc_oh_reg[101][3] + loc_oh_reg[102][3] + loc_oh_reg[103][3] + loc_oh_reg[104][3] + loc_oh_reg[105][3] + loc_oh_reg[106][3] + loc_oh_reg[107][3] + loc_oh_reg[108][3] + loc_oh_reg[109][3] + loc_oh_reg[110][3] + loc_oh_reg[111][3] + loc_oh_reg[112][3] + loc_oh_reg[113][3] + loc_oh_reg[114][3] + loc_oh_reg[115][3] + loc_oh_reg[116][3] + loc_oh_reg[117][3] + loc_oh_reg[118][3] + loc_oh_reg[119][3] + loc_oh_reg[120][3] + loc_oh_reg[121][3] + loc_oh_reg[122][3] + loc_oh_reg[123][3] + loc_oh_reg[124][3] + loc_oh_reg[125][3] + loc_oh_reg[126][3] + loc_oh_reg[127][3];
    n_dsum_reg[28] = loc_oh_reg[128][3] + loc_oh_reg[129][3] + loc_oh_reg[130][3] + loc_oh_reg[131][3] + loc_oh_reg[132][3] + loc_oh_reg[133][3] + loc_oh_reg[134][3] + loc_oh_reg[135][3] + loc_oh_reg[136][3] + loc_oh_reg[137][3] + loc_oh_reg[138][3] + loc_oh_reg[139][3] + loc_oh_reg[140][3] + loc_oh_reg[141][3] + loc_oh_reg[142][3] + loc_oh_reg[143][3] + loc_oh_reg[144][3] + loc_oh_reg[145][3] + loc_oh_reg[146][3] + loc_oh_reg[147][3] + loc_oh_reg[148][3] + loc_oh_reg[149][3] + loc_oh_reg[150][3] + loc_oh_reg[151][3] + loc_oh_reg[152][3] + loc_oh_reg[153][3] + loc_oh_reg[154][3] + loc_oh_reg[155][3] + loc_oh_reg[156][3] + loc_oh_reg[157][3] + loc_oh_reg[158][3] + loc_oh_reg[159][3];
    n_dsum_reg[29] = loc_oh_reg[160][3] + loc_oh_reg[161][3] + loc_oh_reg[162][3] + loc_oh_reg[163][3] + loc_oh_reg[164][3] + loc_oh_reg[165][3] + loc_oh_reg[166][3] + loc_oh_reg[167][3] + loc_oh_reg[168][3] + loc_oh_reg[169][3] + loc_oh_reg[170][3] + loc_oh_reg[171][3] + loc_oh_reg[172][3] + loc_oh_reg[173][3] + loc_oh_reg[174][3] + loc_oh_reg[175][3] + loc_oh_reg[176][3] + loc_oh_reg[177][3] + loc_oh_reg[178][3] + loc_oh_reg[179][3] + loc_oh_reg[180][3] + loc_oh_reg[181][3] + loc_oh_reg[182][3] + loc_oh_reg[183][3] + loc_oh_reg[184][3] + loc_oh_reg[185][3] + loc_oh_reg[186][3] + loc_oh_reg[187][3] + loc_oh_reg[188][3] + loc_oh_reg[189][3] + loc_oh_reg[190][3] + loc_oh_reg[191][3];
    n_dsum_reg[30] = loc_oh_reg[192][3] + loc_oh_reg[193][3] + loc_oh_reg[194][3] + loc_oh_reg[195][3] + loc_oh_reg[196][3] + loc_oh_reg[197][3] + loc_oh_reg[198][3] + loc_oh_reg[199][3] + loc_oh_reg[200][3] + loc_oh_reg[201][3] + loc_oh_reg[202][3] + loc_oh_reg[203][3] + loc_oh_reg[204][3] + loc_oh_reg[205][3] + loc_oh_reg[206][3] + loc_oh_reg[207][3] + loc_oh_reg[208][3] + loc_oh_reg[209][3] + loc_oh_reg[210][3] + loc_oh_reg[211][3] + loc_oh_reg[212][3] + loc_oh_reg[213][3] + loc_oh_reg[214][3] + loc_oh_reg[215][3] + loc_oh_reg[216][3] + loc_oh_reg[217][3] + loc_oh_reg[218][3] + loc_oh_reg[219][3] + loc_oh_reg[220][3] + loc_oh_reg[221][3] + loc_oh_reg[222][3] + loc_oh_reg[223][3];
    n_dsum_reg[31] = loc_oh_reg[224][3] + loc_oh_reg[225][3] + loc_oh_reg[226][3] + loc_oh_reg[227][3] + loc_oh_reg[228][3] + loc_oh_reg[229][3] + loc_oh_reg[230][3] + loc_oh_reg[231][3] + loc_oh_reg[232][3] + loc_oh_reg[233][3] + loc_oh_reg[234][3] + loc_oh_reg[235][3] + loc_oh_reg[236][3] + loc_oh_reg[237][3] + loc_oh_reg[238][3] + loc_oh_reg[239][3] + loc_oh_reg[240][3] + loc_oh_reg[241][3] + loc_oh_reg[242][3] + loc_oh_reg[243][3] + loc_oh_reg[244][3] + loc_oh_reg[245][3] + loc_oh_reg[246][3] + loc_oh_reg[247][3] + loc_oh_reg[248][3] + loc_oh_reg[249][3] + loc_oh_reg[250][3] + loc_oh_reg[251][3] + loc_oh_reg[252][3] + loc_oh_reg[253][3] + loc_oh_reg[254][3] + loc_oh_reg[255][3];

    n_dsum_reg[32] = loc_oh_reg[0][4] + loc_oh_reg[1][4] + loc_oh_reg[2][4] + loc_oh_reg[3][4] + loc_oh_reg[4][4] + loc_oh_reg[5][4] + loc_oh_reg[6][4] + loc_oh_reg[7][4] + loc_oh_reg[8][4] + loc_oh_reg[9][4] + loc_oh_reg[10][4] + loc_oh_reg[11][4] + loc_oh_reg[12][4] + loc_oh_reg[13][4] + loc_oh_reg[14][4] + loc_oh_reg[15][4] + loc_oh_reg[16][4] + loc_oh_reg[17][4] + loc_oh_reg[18][4] + loc_oh_reg[19][4] + loc_oh_reg[20][4] + loc_oh_reg[21][4] + loc_oh_reg[22][4] + loc_oh_reg[23][4] + loc_oh_reg[24][4] + loc_oh_reg[25][4] + loc_oh_reg[26][4] + loc_oh_reg[27][4] + loc_oh_reg[28][4] + loc_oh_reg[29][4] + loc_oh_reg[30][4] + loc_oh_reg[31][4];
    n_dsum_reg[33] = loc_oh_reg[32][4] + loc_oh_reg[33][4] + loc_oh_reg[34][4] + loc_oh_reg[35][4] + loc_oh_reg[36][4] + loc_oh_reg[37][4] + loc_oh_reg[38][4] + loc_oh_reg[39][4] + loc_oh_reg[40][4] + loc_oh_reg[41][4] + loc_oh_reg[42][4] + loc_oh_reg[43][4] + loc_oh_reg[44][4] + loc_oh_reg[45][4] + loc_oh_reg[46][4] + loc_oh_reg[47][4] + loc_oh_reg[48][4] + loc_oh_reg[49][4] + loc_oh_reg[50][4] + loc_oh_reg[51][4] + loc_oh_reg[52][4] + loc_oh_reg[53][4] + loc_oh_reg[54][4] + loc_oh_reg[55][4] + loc_oh_reg[56][4] + loc_oh_reg[57][4] + loc_oh_reg[58][4] + loc_oh_reg[59][4] + loc_oh_reg[60][4] + loc_oh_reg[61][4] + loc_oh_reg[62][4] + loc_oh_reg[63][4];
    n_dsum_reg[34] = loc_oh_reg[64][4] + loc_oh_reg[65][4] + loc_oh_reg[66][4] + loc_oh_reg[67][4] + loc_oh_reg[68][4] + loc_oh_reg[69][4] + loc_oh_reg[70][4] + loc_oh_reg[71][4] + loc_oh_reg[72][4] + loc_oh_reg[73][4] + loc_oh_reg[74][4] + loc_oh_reg[75][4] + loc_oh_reg[76][4] + loc_oh_reg[77][4] + loc_oh_reg[78][4] + loc_oh_reg[79][4] + loc_oh_reg[80][4] + loc_oh_reg[81][4] + loc_oh_reg[82][4] + loc_oh_reg[83][4] + loc_oh_reg[84][4] + loc_oh_reg[85][4] + loc_oh_reg[86][4] + loc_oh_reg[87][4] + loc_oh_reg[88][4] + loc_oh_reg[89][4] + loc_oh_reg[90][4] + loc_oh_reg[91][4] + loc_oh_reg[92][4] + loc_oh_reg[93][4] + loc_oh_reg[94][4] + loc_oh_reg[95][4];
    n_dsum_reg[35] = loc_oh_reg[96][4] + loc_oh_reg[97][4] + loc_oh_reg[98][4] + loc_oh_reg[99][4] + loc_oh_reg[100][4] + loc_oh_reg[101][4] + loc_oh_reg[102][4] + loc_oh_reg[103][4] + loc_oh_reg[104][4] + loc_oh_reg[105][4] + loc_oh_reg[106][4] + loc_oh_reg[107][4] + loc_oh_reg[108][4] + loc_oh_reg[109][4] + loc_oh_reg[110][4] + loc_oh_reg[111][4] + loc_oh_reg[112][4] + loc_oh_reg[113][4] + loc_oh_reg[114][4] + loc_oh_reg[115][4] + loc_oh_reg[116][4] + loc_oh_reg[117][4] + loc_oh_reg[118][4] + loc_oh_reg[119][4] + loc_oh_reg[120][4] + loc_oh_reg[121][4] + loc_oh_reg[122][4] + loc_oh_reg[123][4] + loc_oh_reg[124][4] + loc_oh_reg[125][4] + loc_oh_reg[126][4] + loc_oh_reg[127][4];
    n_dsum_reg[36] = loc_oh_reg[128][4] + loc_oh_reg[129][4] + loc_oh_reg[130][4] + loc_oh_reg[131][4] + loc_oh_reg[132][4] + loc_oh_reg[133][4] + loc_oh_reg[134][4] + loc_oh_reg[135][4] + loc_oh_reg[136][4] + loc_oh_reg[137][4] + loc_oh_reg[138][4] + loc_oh_reg[139][4] + loc_oh_reg[140][4] + loc_oh_reg[141][4] + loc_oh_reg[142][4] + loc_oh_reg[143][4] + loc_oh_reg[144][4] + loc_oh_reg[145][4] + loc_oh_reg[146][4] + loc_oh_reg[147][4] + loc_oh_reg[148][4] + loc_oh_reg[149][4] + loc_oh_reg[150][4] + loc_oh_reg[151][4] + loc_oh_reg[152][4] + loc_oh_reg[153][4] + loc_oh_reg[154][4] + loc_oh_reg[155][4] + loc_oh_reg[156][4] + loc_oh_reg[157][4] + loc_oh_reg[158][4] + loc_oh_reg[159][4];
    n_dsum_reg[37] = loc_oh_reg[160][4] + loc_oh_reg[161][4] + loc_oh_reg[162][4] + loc_oh_reg[163][4] + loc_oh_reg[164][4] + loc_oh_reg[165][4] + loc_oh_reg[166][4] + loc_oh_reg[167][4] + loc_oh_reg[168][4] + loc_oh_reg[169][4] + loc_oh_reg[170][4] + loc_oh_reg[171][4] + loc_oh_reg[172][4] + loc_oh_reg[173][4] + loc_oh_reg[174][4] + loc_oh_reg[175][4] + loc_oh_reg[176][4] + loc_oh_reg[177][4] + loc_oh_reg[178][4] + loc_oh_reg[179][4] + loc_oh_reg[180][4] + loc_oh_reg[181][4] + loc_oh_reg[182][4] + loc_oh_reg[183][4] + loc_oh_reg[184][4] + loc_oh_reg[185][4] + loc_oh_reg[186][4] + loc_oh_reg[187][4] + loc_oh_reg[188][4] + loc_oh_reg[189][4] + loc_oh_reg[190][4] + loc_oh_reg[191][4];
    n_dsum_reg[38] = loc_oh_reg[192][4] + loc_oh_reg[193][4] + loc_oh_reg[194][4] + loc_oh_reg[195][4] + loc_oh_reg[196][4] + loc_oh_reg[197][4] + loc_oh_reg[198][4] + loc_oh_reg[199][4] + loc_oh_reg[200][4] + loc_oh_reg[201][4] + loc_oh_reg[202][4] + loc_oh_reg[203][4] + loc_oh_reg[204][4] + loc_oh_reg[205][4] + loc_oh_reg[206][4] + loc_oh_reg[207][4] + loc_oh_reg[208][4] + loc_oh_reg[209][4] + loc_oh_reg[210][4] + loc_oh_reg[211][4] + loc_oh_reg[212][4] + loc_oh_reg[213][4] + loc_oh_reg[214][4] + loc_oh_reg[215][4] + loc_oh_reg[216][4] + loc_oh_reg[217][4] + loc_oh_reg[218][4] + loc_oh_reg[219][4] + loc_oh_reg[220][4] + loc_oh_reg[221][4] + loc_oh_reg[222][4] + loc_oh_reg[223][4];
    n_dsum_reg[39] = loc_oh_reg[224][4] + loc_oh_reg[225][4] + loc_oh_reg[226][4] + loc_oh_reg[227][4] + loc_oh_reg[228][4] + loc_oh_reg[229][4] + loc_oh_reg[230][4] + loc_oh_reg[231][4] + loc_oh_reg[232][4] + loc_oh_reg[233][4] + loc_oh_reg[234][4] + loc_oh_reg[235][4] + loc_oh_reg[236][4] + loc_oh_reg[237][4] + loc_oh_reg[238][4] + loc_oh_reg[239][4] + loc_oh_reg[240][4] + loc_oh_reg[241][4] + loc_oh_reg[242][4] + loc_oh_reg[243][4] + loc_oh_reg[244][4] + loc_oh_reg[245][4] + loc_oh_reg[246][4] + loc_oh_reg[247][4] + loc_oh_reg[248][4] + loc_oh_reg[249][4] + loc_oh_reg[250][4] + loc_oh_reg[251][4] + loc_oh_reg[252][4] + loc_oh_reg[253][4] + loc_oh_reg[254][4] + loc_oh_reg[255][4];

    n_dsum_reg[40] = loc_oh_reg[0][5] + loc_oh_reg[1][5] + loc_oh_reg[2][5] + loc_oh_reg[3][5] + loc_oh_reg[4][5] + loc_oh_reg[5][5] + loc_oh_reg[6][5] + loc_oh_reg[7][5] + loc_oh_reg[8][5] + loc_oh_reg[9][5] + loc_oh_reg[10][5] + loc_oh_reg[11][5] + loc_oh_reg[12][5] + loc_oh_reg[13][5] + loc_oh_reg[14][5] + loc_oh_reg[15][5] + loc_oh_reg[16][5] + loc_oh_reg[17][5] + loc_oh_reg[18][5] + loc_oh_reg[19][5] + loc_oh_reg[20][5] + loc_oh_reg[21][5] + loc_oh_reg[22][5] + loc_oh_reg[23][5] + loc_oh_reg[24][5] + loc_oh_reg[25][5] + loc_oh_reg[26][5] + loc_oh_reg[27][5] + loc_oh_reg[28][5] + loc_oh_reg[29][5] + loc_oh_reg[30][5] + loc_oh_reg[31][5];
    n_dsum_reg[41] = loc_oh_reg[32][5] + loc_oh_reg[33][5] + loc_oh_reg[34][5] + loc_oh_reg[35][5] + loc_oh_reg[36][5] + loc_oh_reg[37][5] + loc_oh_reg[38][5] + loc_oh_reg[39][5] + loc_oh_reg[40][5] + loc_oh_reg[41][5] + loc_oh_reg[42][5] + loc_oh_reg[43][5] + loc_oh_reg[44][5] + loc_oh_reg[45][5] + loc_oh_reg[46][5] + loc_oh_reg[47][5] + loc_oh_reg[48][5] + loc_oh_reg[49][5] + loc_oh_reg[50][5] + loc_oh_reg[51][5] + loc_oh_reg[52][5] + loc_oh_reg[53][5] + loc_oh_reg[54][5] + loc_oh_reg[55][5] + loc_oh_reg[56][5] + loc_oh_reg[57][5] + loc_oh_reg[58][5] + loc_oh_reg[59][5] + loc_oh_reg[60][5] + loc_oh_reg[61][5] + loc_oh_reg[62][5] + loc_oh_reg[63][5];
    n_dsum_reg[42] = loc_oh_reg[64][5] + loc_oh_reg[65][5] + loc_oh_reg[66][5] + loc_oh_reg[67][5] + loc_oh_reg[68][5] + loc_oh_reg[69][5] + loc_oh_reg[70][5] + loc_oh_reg[71][5] + loc_oh_reg[72][5] + loc_oh_reg[73][5] + loc_oh_reg[74][5] + loc_oh_reg[75][5] + loc_oh_reg[76][5] + loc_oh_reg[77][5] + loc_oh_reg[78][5] + loc_oh_reg[79][5] + loc_oh_reg[80][5] + loc_oh_reg[81][5] + loc_oh_reg[82][5] + loc_oh_reg[83][5] + loc_oh_reg[84][5] + loc_oh_reg[85][5] + loc_oh_reg[86][5] + loc_oh_reg[87][5] + loc_oh_reg[88][5] + loc_oh_reg[89][5] + loc_oh_reg[90][5] + loc_oh_reg[91][5] + loc_oh_reg[92][5] + loc_oh_reg[93][5] + loc_oh_reg[94][5] + loc_oh_reg[95][5];
    n_dsum_reg[43] = loc_oh_reg[96][5] + loc_oh_reg[97][5] + loc_oh_reg[98][5] + loc_oh_reg[99][5] + loc_oh_reg[100][5] + loc_oh_reg[101][5] + loc_oh_reg[102][5] + loc_oh_reg[103][5] + loc_oh_reg[104][5] + loc_oh_reg[105][5] + loc_oh_reg[106][5] + loc_oh_reg[107][5] + loc_oh_reg[108][5] + loc_oh_reg[109][5] + loc_oh_reg[110][5] + loc_oh_reg[111][5] + loc_oh_reg[112][5] + loc_oh_reg[113][5] + loc_oh_reg[114][5] + loc_oh_reg[115][5] + loc_oh_reg[116][5] + loc_oh_reg[117][5] + loc_oh_reg[118][5] + loc_oh_reg[119][5] + loc_oh_reg[120][5] + loc_oh_reg[121][5] + loc_oh_reg[122][5] + loc_oh_reg[123][5] + loc_oh_reg[124][5] + loc_oh_reg[125][5] + loc_oh_reg[126][5] + loc_oh_reg[127][5];
    n_dsum_reg[44] = loc_oh_reg[128][5] + loc_oh_reg[129][5] + loc_oh_reg[130][5] + loc_oh_reg[131][5] + loc_oh_reg[132][5] + loc_oh_reg[133][5] + loc_oh_reg[134][5] + loc_oh_reg[135][5] + loc_oh_reg[136][5] + loc_oh_reg[137][5] + loc_oh_reg[138][5] + loc_oh_reg[139][5] + loc_oh_reg[140][5] + loc_oh_reg[141][5] + loc_oh_reg[142][5] + loc_oh_reg[143][5] + loc_oh_reg[144][5] + loc_oh_reg[145][5] + loc_oh_reg[146][5] + loc_oh_reg[147][5] + loc_oh_reg[148][5] + loc_oh_reg[149][5] + loc_oh_reg[150][5] + loc_oh_reg[151][5] + loc_oh_reg[152][5] + loc_oh_reg[153][5] + loc_oh_reg[154][5] + loc_oh_reg[155][5] + loc_oh_reg[156][5] + loc_oh_reg[157][5] + loc_oh_reg[158][5] + loc_oh_reg[159][5];
    n_dsum_reg[45] = loc_oh_reg[160][5] + loc_oh_reg[161][5] + loc_oh_reg[162][5] + loc_oh_reg[163][5] + loc_oh_reg[164][5] + loc_oh_reg[165][5] + loc_oh_reg[166][5] + loc_oh_reg[167][5] + loc_oh_reg[168][5] + loc_oh_reg[169][5] + loc_oh_reg[170][5] + loc_oh_reg[171][5] + loc_oh_reg[172][5] + loc_oh_reg[173][5] + loc_oh_reg[174][5] + loc_oh_reg[175][5] + loc_oh_reg[176][5] + loc_oh_reg[177][5] + loc_oh_reg[178][5] + loc_oh_reg[179][5] + loc_oh_reg[180][5] + loc_oh_reg[181][5] + loc_oh_reg[182][5] + loc_oh_reg[183][5] + loc_oh_reg[184][5] + loc_oh_reg[185][5] + loc_oh_reg[186][5] + loc_oh_reg[187][5] + loc_oh_reg[188][5] + loc_oh_reg[189][5] + loc_oh_reg[190][5] + loc_oh_reg[191][5];
    n_dsum_reg[46] = loc_oh_reg[192][5] + loc_oh_reg[193][5] + loc_oh_reg[194][5] + loc_oh_reg[195][5] + loc_oh_reg[196][5] + loc_oh_reg[197][5] + loc_oh_reg[198][5] + loc_oh_reg[199][5] + loc_oh_reg[200][5] + loc_oh_reg[201][5] + loc_oh_reg[202][5] + loc_oh_reg[203][5] + loc_oh_reg[204][5] + loc_oh_reg[205][5] + loc_oh_reg[206][5] + loc_oh_reg[207][5] + loc_oh_reg[208][5] + loc_oh_reg[209][5] + loc_oh_reg[210][5] + loc_oh_reg[211][5] + loc_oh_reg[212][5] + loc_oh_reg[213][5] + loc_oh_reg[214][5] + loc_oh_reg[215][5] + loc_oh_reg[216][5] + loc_oh_reg[217][5] + loc_oh_reg[218][5] + loc_oh_reg[219][5] + loc_oh_reg[220][5] + loc_oh_reg[221][5] + loc_oh_reg[222][5] + loc_oh_reg[223][5];
    n_dsum_reg[47] = loc_oh_reg[224][5] + loc_oh_reg[225][5] + loc_oh_reg[226][5] + loc_oh_reg[227][5] + loc_oh_reg[228][5] + loc_oh_reg[229][5] + loc_oh_reg[230][5] + loc_oh_reg[231][5] + loc_oh_reg[232][5] + loc_oh_reg[233][5] + loc_oh_reg[234][5] + loc_oh_reg[235][5] + loc_oh_reg[236][5] + loc_oh_reg[237][5] + loc_oh_reg[238][5] + loc_oh_reg[239][5] + loc_oh_reg[240][5] + loc_oh_reg[241][5] + loc_oh_reg[242][5] + loc_oh_reg[243][5] + loc_oh_reg[244][5] + loc_oh_reg[245][5] + loc_oh_reg[246][5] + loc_oh_reg[247][5] + loc_oh_reg[248][5] + loc_oh_reg[249][5] + loc_oh_reg[250][5] + loc_oh_reg[251][5] + loc_oh_reg[252][5] + loc_oh_reg[253][5] + loc_oh_reg[254][5] + loc_oh_reg[255][5];

    n_dsum_reg[48] = loc_oh_reg[0][6] + loc_oh_reg[1][6] + loc_oh_reg[2][6] + loc_oh_reg[3][6] + loc_oh_reg[4][6] + loc_oh_reg[5][6] + loc_oh_reg[6][6] + loc_oh_reg[7][6] + loc_oh_reg[8][6] + loc_oh_reg[9][6] + loc_oh_reg[10][6] + loc_oh_reg[11][6] + loc_oh_reg[12][6] + loc_oh_reg[13][6] + loc_oh_reg[14][6] + loc_oh_reg[15][6] + loc_oh_reg[16][6] + loc_oh_reg[17][6] + loc_oh_reg[18][6] + loc_oh_reg[19][6] + loc_oh_reg[20][6] + loc_oh_reg[21][6] + loc_oh_reg[22][6] + loc_oh_reg[23][6] + loc_oh_reg[24][6] + loc_oh_reg[25][6] + loc_oh_reg[26][6] + loc_oh_reg[27][6] + loc_oh_reg[28][6] + loc_oh_reg[29][6] + loc_oh_reg[30][6] + loc_oh_reg[31][6];
    n_dsum_reg[49] = loc_oh_reg[32][6] + loc_oh_reg[33][6] + loc_oh_reg[34][6] + loc_oh_reg[35][6] + loc_oh_reg[36][6] + loc_oh_reg[37][6] + loc_oh_reg[38][6] + loc_oh_reg[39][6] + loc_oh_reg[40][6] + loc_oh_reg[41][6] + loc_oh_reg[42][6] + loc_oh_reg[43][6] + loc_oh_reg[44][6] + loc_oh_reg[45][6] + loc_oh_reg[46][6] + loc_oh_reg[47][6] + loc_oh_reg[48][6] + loc_oh_reg[49][6] + loc_oh_reg[50][6] + loc_oh_reg[51][6] + loc_oh_reg[52][6] + loc_oh_reg[53][6] + loc_oh_reg[54][6] + loc_oh_reg[55][6] + loc_oh_reg[56][6] + loc_oh_reg[57][6] + loc_oh_reg[58][6] + loc_oh_reg[59][6] + loc_oh_reg[60][6] + loc_oh_reg[61][6] + loc_oh_reg[62][6] + loc_oh_reg[63][6];
    n_dsum_reg[50] = loc_oh_reg[64][6] + loc_oh_reg[65][6] + loc_oh_reg[66][6] + loc_oh_reg[67][6] + loc_oh_reg[68][6] + loc_oh_reg[69][6] + loc_oh_reg[70][6] + loc_oh_reg[71][6] + loc_oh_reg[72][6] + loc_oh_reg[73][6] + loc_oh_reg[74][6] + loc_oh_reg[75][6] + loc_oh_reg[76][6] + loc_oh_reg[77][6] + loc_oh_reg[78][6] + loc_oh_reg[79][6] + loc_oh_reg[80][6] + loc_oh_reg[81][6] + loc_oh_reg[82][6] + loc_oh_reg[83][6] + loc_oh_reg[84][6] + loc_oh_reg[85][6] + loc_oh_reg[86][6] + loc_oh_reg[87][6] + loc_oh_reg[88][6] + loc_oh_reg[89][6] + loc_oh_reg[90][6] + loc_oh_reg[91][6] + loc_oh_reg[92][6] + loc_oh_reg[93][6] + loc_oh_reg[94][6] + loc_oh_reg[95][6];
    n_dsum_reg[51] = loc_oh_reg[96][6] + loc_oh_reg[97][6] + loc_oh_reg[98][6] + loc_oh_reg[99][6] + loc_oh_reg[100][6] + loc_oh_reg[101][6] + loc_oh_reg[102][6] + loc_oh_reg[103][6] + loc_oh_reg[104][6] + loc_oh_reg[105][6] + loc_oh_reg[106][6] + loc_oh_reg[107][6] + loc_oh_reg[108][6] + loc_oh_reg[109][6] + loc_oh_reg[110][6] + loc_oh_reg[111][6] + loc_oh_reg[112][6] + loc_oh_reg[113][6] + loc_oh_reg[114][6] + loc_oh_reg[115][6] + loc_oh_reg[116][6] + loc_oh_reg[117][6] + loc_oh_reg[118][6] + loc_oh_reg[119][6] + loc_oh_reg[120][6] + loc_oh_reg[121][6] + loc_oh_reg[122][6] + loc_oh_reg[123][6] + loc_oh_reg[124][6] + loc_oh_reg[125][6] + loc_oh_reg[126][6] + loc_oh_reg[127][6];
    n_dsum_reg[52] = loc_oh_reg[128][6] + loc_oh_reg[129][6] + loc_oh_reg[130][6] + loc_oh_reg[131][6] + loc_oh_reg[132][6] + loc_oh_reg[133][6] + loc_oh_reg[134][6] + loc_oh_reg[135][6] + loc_oh_reg[136][6] + loc_oh_reg[137][6] + loc_oh_reg[138][6] + loc_oh_reg[139][6] + loc_oh_reg[140][6] + loc_oh_reg[141][6] + loc_oh_reg[142][6] + loc_oh_reg[143][6] + loc_oh_reg[144][6] + loc_oh_reg[145][6] + loc_oh_reg[146][6] + loc_oh_reg[147][6] + loc_oh_reg[148][6] + loc_oh_reg[149][6] + loc_oh_reg[150][6] + loc_oh_reg[151][6] + loc_oh_reg[152][6] + loc_oh_reg[153][6] + loc_oh_reg[154][6] + loc_oh_reg[155][6] + loc_oh_reg[156][6] + loc_oh_reg[157][6] + loc_oh_reg[158][6] + loc_oh_reg[159][6];
    n_dsum_reg[53] = loc_oh_reg[160][6] + loc_oh_reg[161][6] + loc_oh_reg[162][6] + loc_oh_reg[163][6] + loc_oh_reg[164][6] + loc_oh_reg[165][6] + loc_oh_reg[166][6] + loc_oh_reg[167][6] + loc_oh_reg[168][6] + loc_oh_reg[169][6] + loc_oh_reg[170][6] + loc_oh_reg[171][6] + loc_oh_reg[172][6] + loc_oh_reg[173][6] + loc_oh_reg[174][6] + loc_oh_reg[175][6] + loc_oh_reg[176][6] + loc_oh_reg[177][6] + loc_oh_reg[178][6] + loc_oh_reg[179][6] + loc_oh_reg[180][6] + loc_oh_reg[181][6] + loc_oh_reg[182][6] + loc_oh_reg[183][6] + loc_oh_reg[184][6] + loc_oh_reg[185][6] + loc_oh_reg[186][6] + loc_oh_reg[187][6] + loc_oh_reg[188][6] + loc_oh_reg[189][6] + loc_oh_reg[190][6] + loc_oh_reg[191][6];
    n_dsum_reg[54] = loc_oh_reg[192][6] + loc_oh_reg[193][6] + loc_oh_reg[194][6] + loc_oh_reg[195][6] + loc_oh_reg[196][6] + loc_oh_reg[197][6] + loc_oh_reg[198][6] + loc_oh_reg[199][6] + loc_oh_reg[200][6] + loc_oh_reg[201][6] + loc_oh_reg[202][6] + loc_oh_reg[203][6] + loc_oh_reg[204][6] + loc_oh_reg[205][6] + loc_oh_reg[206][6] + loc_oh_reg[207][6] + loc_oh_reg[208][6] + loc_oh_reg[209][6] + loc_oh_reg[210][6] + loc_oh_reg[211][6] + loc_oh_reg[212][6] + loc_oh_reg[213][6] + loc_oh_reg[214][6] + loc_oh_reg[215][6] + loc_oh_reg[216][6] + loc_oh_reg[217][6] + loc_oh_reg[218][6] + loc_oh_reg[219][6] + loc_oh_reg[220][6] + loc_oh_reg[221][6] + loc_oh_reg[222][6] + loc_oh_reg[223][6];
    n_dsum_reg[55] = loc_oh_reg[224][6] + loc_oh_reg[225][6] + loc_oh_reg[226][6] + loc_oh_reg[227][6] + loc_oh_reg[228][6] + loc_oh_reg[229][6] + loc_oh_reg[230][6] + loc_oh_reg[231][6] + loc_oh_reg[232][6] + loc_oh_reg[233][6] + loc_oh_reg[234][6] + loc_oh_reg[235][6] + loc_oh_reg[236][6] + loc_oh_reg[237][6] + loc_oh_reg[238][6] + loc_oh_reg[239][6] + loc_oh_reg[240][6] + loc_oh_reg[241][6] + loc_oh_reg[242][6] + loc_oh_reg[243][6] + loc_oh_reg[244][6] + loc_oh_reg[245][6] + loc_oh_reg[246][6] + loc_oh_reg[247][6] + loc_oh_reg[248][6] + loc_oh_reg[249][6] + loc_oh_reg[250][6] + loc_oh_reg[251][6] + loc_oh_reg[252][6] + loc_oh_reg[253][6] + loc_oh_reg[254][6] + loc_oh_reg[255][6];

    n_dsum_reg[56] = loc_oh_reg[0][7] + loc_oh_reg[1][7] + loc_oh_reg[2][7] + loc_oh_reg[3][7] + loc_oh_reg[4][7] + loc_oh_reg[5][7] + loc_oh_reg[6][7] + loc_oh_reg[7][7] + loc_oh_reg[8][7] + loc_oh_reg[9][7] + loc_oh_reg[10][7] + loc_oh_reg[11][7] + loc_oh_reg[12][7] + loc_oh_reg[13][7] + loc_oh_reg[14][7] + loc_oh_reg[15][7] + loc_oh_reg[16][7] + loc_oh_reg[17][7] + loc_oh_reg[18][7] + loc_oh_reg[19][7] + loc_oh_reg[20][7] + loc_oh_reg[21][7] + loc_oh_reg[22][7] + loc_oh_reg[23][7] + loc_oh_reg[24][7] + loc_oh_reg[25][7] + loc_oh_reg[26][7] + loc_oh_reg[27][7] + loc_oh_reg[28][7] + loc_oh_reg[29][7] + loc_oh_reg[30][7] + loc_oh_reg[31][7];
    n_dsum_reg[57] = loc_oh_reg[32][7] + loc_oh_reg[33][7] + loc_oh_reg[34][7] + loc_oh_reg[35][7] + loc_oh_reg[36][7] + loc_oh_reg[37][7] + loc_oh_reg[38][7] + loc_oh_reg[39][7] + loc_oh_reg[40][7] + loc_oh_reg[41][7] + loc_oh_reg[42][7] + loc_oh_reg[43][7] + loc_oh_reg[44][7] + loc_oh_reg[45][7] + loc_oh_reg[46][7] + loc_oh_reg[47][7] + loc_oh_reg[48][7] + loc_oh_reg[49][7] + loc_oh_reg[50][7] + loc_oh_reg[51][7] + loc_oh_reg[52][7] + loc_oh_reg[53][7] + loc_oh_reg[54][7] + loc_oh_reg[55][7] + loc_oh_reg[56][7] + loc_oh_reg[57][7] + loc_oh_reg[58][7] + loc_oh_reg[59][7] + loc_oh_reg[60][7] + loc_oh_reg[61][7] + loc_oh_reg[62][7] + loc_oh_reg[63][7];
    n_dsum_reg[58] = loc_oh_reg[64][7] + loc_oh_reg[65][7] + loc_oh_reg[66][7] + loc_oh_reg[67][7] + loc_oh_reg[68][7] + loc_oh_reg[69][7] + loc_oh_reg[70][7] + loc_oh_reg[71][7] + loc_oh_reg[72][7] + loc_oh_reg[73][7] + loc_oh_reg[74][7] + loc_oh_reg[75][7] + loc_oh_reg[76][7] + loc_oh_reg[77][7] + loc_oh_reg[78][7] + loc_oh_reg[79][7] + loc_oh_reg[80][7] + loc_oh_reg[81][7] + loc_oh_reg[82][7] + loc_oh_reg[83][7] + loc_oh_reg[84][7] + loc_oh_reg[85][7] + loc_oh_reg[86][7] + loc_oh_reg[87][7] + loc_oh_reg[88][7] + loc_oh_reg[89][7] + loc_oh_reg[90][7] + loc_oh_reg[91][7] + loc_oh_reg[92][7] + loc_oh_reg[93][7] + loc_oh_reg[94][7] + loc_oh_reg[95][7];
    n_dsum_reg[59] = loc_oh_reg[96][7] + loc_oh_reg[97][7] + loc_oh_reg[98][7] + loc_oh_reg[99][7] + loc_oh_reg[100][7] + loc_oh_reg[101][7] + loc_oh_reg[102][7] + loc_oh_reg[103][7] + loc_oh_reg[104][7] + loc_oh_reg[105][7] + loc_oh_reg[106][7] + loc_oh_reg[107][7] + loc_oh_reg[108][7] + loc_oh_reg[109][7] + loc_oh_reg[110][7] + loc_oh_reg[111][7] + loc_oh_reg[112][7] + loc_oh_reg[113][7] + loc_oh_reg[114][7] + loc_oh_reg[115][7] + loc_oh_reg[116][7] + loc_oh_reg[117][7] + loc_oh_reg[118][7] + loc_oh_reg[119][7] + loc_oh_reg[120][7] + loc_oh_reg[121][7] + loc_oh_reg[122][7] + loc_oh_reg[123][7] + loc_oh_reg[124][7] + loc_oh_reg[125][7] + loc_oh_reg[126][7] + loc_oh_reg[127][7];
    n_dsum_reg[60] = loc_oh_reg[128][7] + loc_oh_reg[129][7] + loc_oh_reg[130][7] + loc_oh_reg[131][7] + loc_oh_reg[132][7] + loc_oh_reg[133][7] + loc_oh_reg[134][7] + loc_oh_reg[135][7] + loc_oh_reg[136][7] + loc_oh_reg[137][7] + loc_oh_reg[138][7] + loc_oh_reg[139][7] + loc_oh_reg[140][7] + loc_oh_reg[141][7] + loc_oh_reg[142][7] + loc_oh_reg[143][7] + loc_oh_reg[144][7] + loc_oh_reg[145][7] + loc_oh_reg[146][7] + loc_oh_reg[147][7] + loc_oh_reg[148][7] + loc_oh_reg[149][7] + loc_oh_reg[150][7] + loc_oh_reg[151][7] + loc_oh_reg[152][7] + loc_oh_reg[153][7] + loc_oh_reg[154][7] + loc_oh_reg[155][7] + loc_oh_reg[156][7] + loc_oh_reg[157][7] + loc_oh_reg[158][7] + loc_oh_reg[159][7];
    n_dsum_reg[61] = loc_oh_reg[160][7] + loc_oh_reg[161][7] + loc_oh_reg[162][7] + loc_oh_reg[163][7] + loc_oh_reg[164][7] + loc_oh_reg[165][7] + loc_oh_reg[166][7] + loc_oh_reg[167][7] + loc_oh_reg[168][7] + loc_oh_reg[169][7] + loc_oh_reg[170][7] + loc_oh_reg[171][7] + loc_oh_reg[172][7] + loc_oh_reg[173][7] + loc_oh_reg[174][7] + loc_oh_reg[175][7] + loc_oh_reg[176][7] + loc_oh_reg[177][7] + loc_oh_reg[178][7] + loc_oh_reg[179][7] + loc_oh_reg[180][7] + loc_oh_reg[181][7] + loc_oh_reg[182][7] + loc_oh_reg[183][7] + loc_oh_reg[184][7] + loc_oh_reg[185][7] + loc_oh_reg[186][7] + loc_oh_reg[187][7] + loc_oh_reg[188][7] + loc_oh_reg[189][7] + loc_oh_reg[190][7] + loc_oh_reg[191][7];
    n_dsum_reg[62] = loc_oh_reg[192][7] + loc_oh_reg[193][7] + loc_oh_reg[194][7] + loc_oh_reg[195][7] + loc_oh_reg[196][7] + loc_oh_reg[197][7] + loc_oh_reg[198][7] + loc_oh_reg[199][7] + loc_oh_reg[200][7] + loc_oh_reg[201][7] + loc_oh_reg[202][7] + loc_oh_reg[203][7] + loc_oh_reg[204][7] + loc_oh_reg[205][7] + loc_oh_reg[206][7] + loc_oh_reg[207][7] + loc_oh_reg[208][7] + loc_oh_reg[209][7] + loc_oh_reg[210][7] + loc_oh_reg[211][7] + loc_oh_reg[212][7] + loc_oh_reg[213][7] + loc_oh_reg[214][7] + loc_oh_reg[215][7] + loc_oh_reg[216][7] + loc_oh_reg[217][7] + loc_oh_reg[218][7] + loc_oh_reg[219][7] + loc_oh_reg[220][7] + loc_oh_reg[221][7] + loc_oh_reg[222][7] + loc_oh_reg[223][7];
    n_dsum_reg[63] = loc_oh_reg[224][7] + loc_oh_reg[225][7] + loc_oh_reg[226][7] + loc_oh_reg[227][7] + loc_oh_reg[228][7] + loc_oh_reg[229][7] + loc_oh_reg[230][7] + loc_oh_reg[231][7] + loc_oh_reg[232][7] + loc_oh_reg[233][7] + loc_oh_reg[234][7] + loc_oh_reg[235][7] + loc_oh_reg[236][7] + loc_oh_reg[237][7] + loc_oh_reg[238][7] + loc_oh_reg[239][7] + loc_oh_reg[240][7] + loc_oh_reg[241][7] + loc_oh_reg[242][7] + loc_oh_reg[243][7] + loc_oh_reg[244][7] + loc_oh_reg[245][7] + loc_oh_reg[246][7] + loc_oh_reg[247][7] + loc_oh_reg[248][7] + loc_oh_reg[249][7] + loc_oh_reg[250][7] + loc_oh_reg[251][7] + loc_oh_reg[252][7] + loc_oh_reg[253][7] + loc_oh_reg[254][7] + loc_oh_reg[255][7];

    n_dsum_reg[64] = loc_oh_reg[0][8] + loc_oh_reg[1][8] + loc_oh_reg[2][8] + loc_oh_reg[3][8] + loc_oh_reg[4][8] + loc_oh_reg[5][8] + loc_oh_reg[6][8] + loc_oh_reg[7][8] + loc_oh_reg[8][8] + loc_oh_reg[9][8] + loc_oh_reg[10][8] + loc_oh_reg[11][8] + loc_oh_reg[12][8] + loc_oh_reg[13][8] + loc_oh_reg[14][8] + loc_oh_reg[15][8] + loc_oh_reg[16][8] + loc_oh_reg[17][8] + loc_oh_reg[18][8] + loc_oh_reg[19][8] + loc_oh_reg[20][8] + loc_oh_reg[21][8] + loc_oh_reg[22][8] + loc_oh_reg[23][8] + loc_oh_reg[24][8] + loc_oh_reg[25][8] + loc_oh_reg[26][8] + loc_oh_reg[27][8] + loc_oh_reg[28][8] + loc_oh_reg[29][8] + loc_oh_reg[30][8] + loc_oh_reg[31][8];
    n_dsum_reg[65] = loc_oh_reg[32][8] + loc_oh_reg[33][8] + loc_oh_reg[34][8] + loc_oh_reg[35][8] + loc_oh_reg[36][8] + loc_oh_reg[37][8] + loc_oh_reg[38][8] + loc_oh_reg[39][8] + loc_oh_reg[40][8] + loc_oh_reg[41][8] + loc_oh_reg[42][8] + loc_oh_reg[43][8] + loc_oh_reg[44][8] + loc_oh_reg[45][8] + loc_oh_reg[46][8] + loc_oh_reg[47][8] + loc_oh_reg[48][8] + loc_oh_reg[49][8] + loc_oh_reg[50][8] + loc_oh_reg[51][8] + loc_oh_reg[52][8] + loc_oh_reg[53][8] + loc_oh_reg[54][8] + loc_oh_reg[55][8] + loc_oh_reg[56][8] + loc_oh_reg[57][8] + loc_oh_reg[58][8] + loc_oh_reg[59][8] + loc_oh_reg[60][8] + loc_oh_reg[61][8] + loc_oh_reg[62][8] + loc_oh_reg[63][8];
    n_dsum_reg[66] = loc_oh_reg[64][8] + loc_oh_reg[65][8] + loc_oh_reg[66][8] + loc_oh_reg[67][8] + loc_oh_reg[68][8] + loc_oh_reg[69][8] + loc_oh_reg[70][8] + loc_oh_reg[71][8] + loc_oh_reg[72][8] + loc_oh_reg[73][8] + loc_oh_reg[74][8] + loc_oh_reg[75][8] + loc_oh_reg[76][8] + loc_oh_reg[77][8] + loc_oh_reg[78][8] + loc_oh_reg[79][8] + loc_oh_reg[80][8] + loc_oh_reg[81][8] + loc_oh_reg[82][8] + loc_oh_reg[83][8] + loc_oh_reg[84][8] + loc_oh_reg[85][8] + loc_oh_reg[86][8] + loc_oh_reg[87][8] + loc_oh_reg[88][8] + loc_oh_reg[89][8] + loc_oh_reg[90][8] + loc_oh_reg[91][8] + loc_oh_reg[92][8] + loc_oh_reg[93][8] + loc_oh_reg[94][8] + loc_oh_reg[95][8];
    n_dsum_reg[67] = loc_oh_reg[96][8] + loc_oh_reg[97][8] + loc_oh_reg[98][8] + loc_oh_reg[99][8] + loc_oh_reg[100][8] + loc_oh_reg[101][8] + loc_oh_reg[102][8] + loc_oh_reg[103][8] + loc_oh_reg[104][8] + loc_oh_reg[105][8] + loc_oh_reg[106][8] + loc_oh_reg[107][8] + loc_oh_reg[108][8] + loc_oh_reg[109][8] + loc_oh_reg[110][8] + loc_oh_reg[111][8] + loc_oh_reg[112][8] + loc_oh_reg[113][8] + loc_oh_reg[114][8] + loc_oh_reg[115][8] + loc_oh_reg[116][8] + loc_oh_reg[117][8] + loc_oh_reg[118][8] + loc_oh_reg[119][8] + loc_oh_reg[120][8] + loc_oh_reg[121][8] + loc_oh_reg[122][8] + loc_oh_reg[123][8] + loc_oh_reg[124][8] + loc_oh_reg[125][8] + loc_oh_reg[126][8] + loc_oh_reg[127][8];
    n_dsum_reg[68] = loc_oh_reg[128][8] + loc_oh_reg[129][8] + loc_oh_reg[130][8] + loc_oh_reg[131][8] + loc_oh_reg[132][8] + loc_oh_reg[133][8] + loc_oh_reg[134][8] + loc_oh_reg[135][8] + loc_oh_reg[136][8] + loc_oh_reg[137][8] + loc_oh_reg[138][8] + loc_oh_reg[139][8] + loc_oh_reg[140][8] + loc_oh_reg[141][8] + loc_oh_reg[142][8] + loc_oh_reg[143][8] + loc_oh_reg[144][8] + loc_oh_reg[145][8] + loc_oh_reg[146][8] + loc_oh_reg[147][8] + loc_oh_reg[148][8] + loc_oh_reg[149][8] + loc_oh_reg[150][8] + loc_oh_reg[151][8] + loc_oh_reg[152][8] + loc_oh_reg[153][8] + loc_oh_reg[154][8] + loc_oh_reg[155][8] + loc_oh_reg[156][8] + loc_oh_reg[157][8] + loc_oh_reg[158][8] + loc_oh_reg[159][8];
    n_dsum_reg[69] = loc_oh_reg[160][8] + loc_oh_reg[161][8] + loc_oh_reg[162][8] + loc_oh_reg[163][8] + loc_oh_reg[164][8] + loc_oh_reg[165][8] + loc_oh_reg[166][8] + loc_oh_reg[167][8] + loc_oh_reg[168][8] + loc_oh_reg[169][8] + loc_oh_reg[170][8] + loc_oh_reg[171][8] + loc_oh_reg[172][8] + loc_oh_reg[173][8] + loc_oh_reg[174][8] + loc_oh_reg[175][8] + loc_oh_reg[176][8] + loc_oh_reg[177][8] + loc_oh_reg[178][8] + loc_oh_reg[179][8] + loc_oh_reg[180][8] + loc_oh_reg[181][8] + loc_oh_reg[182][8] + loc_oh_reg[183][8] + loc_oh_reg[184][8] + loc_oh_reg[185][8] + loc_oh_reg[186][8] + loc_oh_reg[187][8] + loc_oh_reg[188][8] + loc_oh_reg[189][8] + loc_oh_reg[190][8] + loc_oh_reg[191][8];
    n_dsum_reg[70] = loc_oh_reg[192][8] + loc_oh_reg[193][8] + loc_oh_reg[194][8] + loc_oh_reg[195][8] + loc_oh_reg[196][8] + loc_oh_reg[197][8] + loc_oh_reg[198][8] + loc_oh_reg[199][8] + loc_oh_reg[200][8] + loc_oh_reg[201][8] + loc_oh_reg[202][8] + loc_oh_reg[203][8] + loc_oh_reg[204][8] + loc_oh_reg[205][8] + loc_oh_reg[206][8] + loc_oh_reg[207][8] + loc_oh_reg[208][8] + loc_oh_reg[209][8] + loc_oh_reg[210][8] + loc_oh_reg[211][8] + loc_oh_reg[212][8] + loc_oh_reg[213][8] + loc_oh_reg[214][8] + loc_oh_reg[215][8] + loc_oh_reg[216][8] + loc_oh_reg[217][8] + loc_oh_reg[218][8] + loc_oh_reg[219][8] + loc_oh_reg[220][8] + loc_oh_reg[221][8] + loc_oh_reg[222][8] + loc_oh_reg[223][8];
    n_dsum_reg[71] = loc_oh_reg[224][8] + loc_oh_reg[225][8] + loc_oh_reg[226][8] + loc_oh_reg[227][8] + loc_oh_reg[228][8] + loc_oh_reg[229][8] + loc_oh_reg[230][8] + loc_oh_reg[231][8] + loc_oh_reg[232][8] + loc_oh_reg[233][8] + loc_oh_reg[234][8] + loc_oh_reg[235][8] + loc_oh_reg[236][8] + loc_oh_reg[237][8] + loc_oh_reg[238][8] + loc_oh_reg[239][8] + loc_oh_reg[240][8] + loc_oh_reg[241][8] + loc_oh_reg[242][8] + loc_oh_reg[243][8] + loc_oh_reg[244][8] + loc_oh_reg[245][8] + loc_oh_reg[246][8] + loc_oh_reg[247][8] + loc_oh_reg[248][8] + loc_oh_reg[249][8] + loc_oh_reg[250][8] + loc_oh_reg[251][8] + loc_oh_reg[252][8] + loc_oh_reg[253][8] + loc_oh_reg[254][8] + loc_oh_reg[255][8];

    n_dsum_reg[72] = loc_oh_reg[0][9] + loc_oh_reg[1][9] + loc_oh_reg[2][9] + loc_oh_reg[3][9] + loc_oh_reg[4][9] + loc_oh_reg[5][9] + loc_oh_reg[6][9] + loc_oh_reg[7][9] + loc_oh_reg[8][9] + loc_oh_reg[9][9] + loc_oh_reg[10][9] + loc_oh_reg[11][9] + loc_oh_reg[12][9] + loc_oh_reg[13][9] + loc_oh_reg[14][9] + loc_oh_reg[15][9] + loc_oh_reg[16][9] + loc_oh_reg[17][9] + loc_oh_reg[18][9] + loc_oh_reg[19][9] + loc_oh_reg[20][9] + loc_oh_reg[21][9] + loc_oh_reg[22][9] + loc_oh_reg[23][9] + loc_oh_reg[24][9] + loc_oh_reg[25][9] + loc_oh_reg[26][9] + loc_oh_reg[27][9] + loc_oh_reg[28][9] + loc_oh_reg[29][9] + loc_oh_reg[30][9] + loc_oh_reg[31][9];
    n_dsum_reg[73] = loc_oh_reg[32][9] + loc_oh_reg[33][9] + loc_oh_reg[34][9] + loc_oh_reg[35][9] + loc_oh_reg[36][9] + loc_oh_reg[37][9] + loc_oh_reg[38][9] + loc_oh_reg[39][9] + loc_oh_reg[40][9] + loc_oh_reg[41][9] + loc_oh_reg[42][9] + loc_oh_reg[43][9] + loc_oh_reg[44][9] + loc_oh_reg[45][9] + loc_oh_reg[46][9] + loc_oh_reg[47][9] + loc_oh_reg[48][9] + loc_oh_reg[49][9] + loc_oh_reg[50][9] + loc_oh_reg[51][9] + loc_oh_reg[52][9] + loc_oh_reg[53][9] + loc_oh_reg[54][9] + loc_oh_reg[55][9] + loc_oh_reg[56][9] + loc_oh_reg[57][9] + loc_oh_reg[58][9] + loc_oh_reg[59][9] + loc_oh_reg[60][9] + loc_oh_reg[61][9] + loc_oh_reg[62][9] + loc_oh_reg[63][9];
    n_dsum_reg[74] = loc_oh_reg[64][9] + loc_oh_reg[65][9] + loc_oh_reg[66][9] + loc_oh_reg[67][9] + loc_oh_reg[68][9] + loc_oh_reg[69][9] + loc_oh_reg[70][9] + loc_oh_reg[71][9] + loc_oh_reg[72][9] + loc_oh_reg[73][9] + loc_oh_reg[74][9] + loc_oh_reg[75][9] + loc_oh_reg[76][9] + loc_oh_reg[77][9] + loc_oh_reg[78][9] + loc_oh_reg[79][9] + loc_oh_reg[80][9] + loc_oh_reg[81][9] + loc_oh_reg[82][9] + loc_oh_reg[83][9] + loc_oh_reg[84][9] + loc_oh_reg[85][9] + loc_oh_reg[86][9] + loc_oh_reg[87][9] + loc_oh_reg[88][9] + loc_oh_reg[89][9] + loc_oh_reg[90][9] + loc_oh_reg[91][9] + loc_oh_reg[92][9] + loc_oh_reg[93][9] + loc_oh_reg[94][9] + loc_oh_reg[95][9];
    n_dsum_reg[75] = loc_oh_reg[96][9] + loc_oh_reg[97][9] + loc_oh_reg[98][9] + loc_oh_reg[99][9] + loc_oh_reg[100][9] + loc_oh_reg[101][9] + loc_oh_reg[102][9] + loc_oh_reg[103][9] + loc_oh_reg[104][9] + loc_oh_reg[105][9] + loc_oh_reg[106][9] + loc_oh_reg[107][9] + loc_oh_reg[108][9] + loc_oh_reg[109][9] + loc_oh_reg[110][9] + loc_oh_reg[111][9] + loc_oh_reg[112][9] + loc_oh_reg[113][9] + loc_oh_reg[114][9] + loc_oh_reg[115][9] + loc_oh_reg[116][9] + loc_oh_reg[117][9] + loc_oh_reg[118][9] + loc_oh_reg[119][9] + loc_oh_reg[120][9] + loc_oh_reg[121][9] + loc_oh_reg[122][9] + loc_oh_reg[123][9] + loc_oh_reg[124][9] + loc_oh_reg[125][9] + loc_oh_reg[126][9] + loc_oh_reg[127][9];
    n_dsum_reg[76] = loc_oh_reg[128][9] + loc_oh_reg[129][9] + loc_oh_reg[130][9] + loc_oh_reg[131][9] + loc_oh_reg[132][9] + loc_oh_reg[133][9] + loc_oh_reg[134][9] + loc_oh_reg[135][9] + loc_oh_reg[136][9] + loc_oh_reg[137][9] + loc_oh_reg[138][9] + loc_oh_reg[139][9] + loc_oh_reg[140][9] + loc_oh_reg[141][9] + loc_oh_reg[142][9] + loc_oh_reg[143][9] + loc_oh_reg[144][9] + loc_oh_reg[145][9] + loc_oh_reg[146][9] + loc_oh_reg[147][9] + loc_oh_reg[148][9] + loc_oh_reg[149][9] + loc_oh_reg[150][9] + loc_oh_reg[151][9] + loc_oh_reg[152][9] + loc_oh_reg[153][9] + loc_oh_reg[154][9] + loc_oh_reg[155][9] + loc_oh_reg[156][9] + loc_oh_reg[157][9] + loc_oh_reg[158][9] + loc_oh_reg[159][9];
    n_dsum_reg[77] = loc_oh_reg[160][9] + loc_oh_reg[161][9] + loc_oh_reg[162][9] + loc_oh_reg[163][9] + loc_oh_reg[164][9] + loc_oh_reg[165][9] + loc_oh_reg[166][9] + loc_oh_reg[167][9] + loc_oh_reg[168][9] + loc_oh_reg[169][9] + loc_oh_reg[170][9] + loc_oh_reg[171][9] + loc_oh_reg[172][9] + loc_oh_reg[173][9] + loc_oh_reg[174][9] + loc_oh_reg[175][9] + loc_oh_reg[176][9] + loc_oh_reg[177][9] + loc_oh_reg[178][9] + loc_oh_reg[179][9] + loc_oh_reg[180][9] + loc_oh_reg[181][9] + loc_oh_reg[182][9] + loc_oh_reg[183][9] + loc_oh_reg[184][9] + loc_oh_reg[185][9] + loc_oh_reg[186][9] + loc_oh_reg[187][9] + loc_oh_reg[188][9] + loc_oh_reg[189][9] + loc_oh_reg[190][9] + loc_oh_reg[191][9];
    n_dsum_reg[78] = loc_oh_reg[192][9] + loc_oh_reg[193][9] + loc_oh_reg[194][9] + loc_oh_reg[195][9] + loc_oh_reg[196][9] + loc_oh_reg[197][9] + loc_oh_reg[198][9] + loc_oh_reg[199][9] + loc_oh_reg[200][9] + loc_oh_reg[201][9] + loc_oh_reg[202][9] + loc_oh_reg[203][9] + loc_oh_reg[204][9] + loc_oh_reg[205][9] + loc_oh_reg[206][9] + loc_oh_reg[207][9] + loc_oh_reg[208][9] + loc_oh_reg[209][9] + loc_oh_reg[210][9] + loc_oh_reg[211][9] + loc_oh_reg[212][9] + loc_oh_reg[213][9] + loc_oh_reg[214][9] + loc_oh_reg[215][9] + loc_oh_reg[216][9] + loc_oh_reg[217][9] + loc_oh_reg[218][9] + loc_oh_reg[219][9] + loc_oh_reg[220][9] + loc_oh_reg[221][9] + loc_oh_reg[222][9] + loc_oh_reg[223][9];
    n_dsum_reg[79] = loc_oh_reg[224][9] + loc_oh_reg[225][9] + loc_oh_reg[226][9] + loc_oh_reg[227][9] + loc_oh_reg[228][9] + loc_oh_reg[229][9] + loc_oh_reg[230][9] + loc_oh_reg[231][9] + loc_oh_reg[232][9] + loc_oh_reg[233][9] + loc_oh_reg[234][9] + loc_oh_reg[235][9] + loc_oh_reg[236][9] + loc_oh_reg[237][9] + loc_oh_reg[238][9] + loc_oh_reg[239][9] + loc_oh_reg[240][9] + loc_oh_reg[241][9] + loc_oh_reg[242][9] + loc_oh_reg[243][9] + loc_oh_reg[244][9] + loc_oh_reg[245][9] + loc_oh_reg[246][9] + loc_oh_reg[247][9] + loc_oh_reg[248][9] + loc_oh_reg[249][9] + loc_oh_reg[250][9] + loc_oh_reg[251][9] + loc_oh_reg[252][9] + loc_oh_reg[253][9] + loc_oh_reg[254][9] + loc_oh_reg[255][9];

    n_dsum_reg[80] = loc_oh_reg[0][10] + loc_oh_reg[1][10] + loc_oh_reg[2][10] + loc_oh_reg[3][10] + loc_oh_reg[4][10] + loc_oh_reg[5][10] + loc_oh_reg[6][10] + loc_oh_reg[7][10] + loc_oh_reg[8][10] + loc_oh_reg[9][10] + loc_oh_reg[10][10] + loc_oh_reg[11][10] + loc_oh_reg[12][10] + loc_oh_reg[13][10] + loc_oh_reg[14][10] + loc_oh_reg[15][10] + loc_oh_reg[16][10] + loc_oh_reg[17][10] + loc_oh_reg[18][10] + loc_oh_reg[19][10] + loc_oh_reg[20][10] + loc_oh_reg[21][10] + loc_oh_reg[22][10] + loc_oh_reg[23][10] + loc_oh_reg[24][10] + loc_oh_reg[25][10] + loc_oh_reg[26][10] + loc_oh_reg[27][10] + loc_oh_reg[28][10] + loc_oh_reg[29][10] + loc_oh_reg[30][10] + loc_oh_reg[31][10];
    n_dsum_reg[81] = loc_oh_reg[32][10] + loc_oh_reg[33][10] + loc_oh_reg[34][10] + loc_oh_reg[35][10] + loc_oh_reg[36][10] + loc_oh_reg[37][10] + loc_oh_reg[38][10] + loc_oh_reg[39][10] + loc_oh_reg[40][10] + loc_oh_reg[41][10] + loc_oh_reg[42][10] + loc_oh_reg[43][10] + loc_oh_reg[44][10] + loc_oh_reg[45][10] + loc_oh_reg[46][10] + loc_oh_reg[47][10] + loc_oh_reg[48][10] + loc_oh_reg[49][10] + loc_oh_reg[50][10] + loc_oh_reg[51][10] + loc_oh_reg[52][10] + loc_oh_reg[53][10] + loc_oh_reg[54][10] + loc_oh_reg[55][10] + loc_oh_reg[56][10] + loc_oh_reg[57][10] + loc_oh_reg[58][10] + loc_oh_reg[59][10] + loc_oh_reg[60][10] + loc_oh_reg[61][10] + loc_oh_reg[62][10] + loc_oh_reg[63][10];
    n_dsum_reg[82] = loc_oh_reg[64][10] + loc_oh_reg[65][10] + loc_oh_reg[66][10] + loc_oh_reg[67][10] + loc_oh_reg[68][10] + loc_oh_reg[69][10] + loc_oh_reg[70][10] + loc_oh_reg[71][10] + loc_oh_reg[72][10] + loc_oh_reg[73][10] + loc_oh_reg[74][10] + loc_oh_reg[75][10] + loc_oh_reg[76][10] + loc_oh_reg[77][10] + loc_oh_reg[78][10] + loc_oh_reg[79][10] + loc_oh_reg[80][10] + loc_oh_reg[81][10] + loc_oh_reg[82][10] + loc_oh_reg[83][10] + loc_oh_reg[84][10] + loc_oh_reg[85][10] + loc_oh_reg[86][10] + loc_oh_reg[87][10] + loc_oh_reg[88][10] + loc_oh_reg[89][10] + loc_oh_reg[90][10] + loc_oh_reg[91][10] + loc_oh_reg[92][10] + loc_oh_reg[93][10] + loc_oh_reg[94][10] + loc_oh_reg[95][10];
    n_dsum_reg[83] = loc_oh_reg[96][10] + loc_oh_reg[97][10] + loc_oh_reg[98][10] + loc_oh_reg[99][10] + loc_oh_reg[100][10] + loc_oh_reg[101][10] + loc_oh_reg[102][10] + loc_oh_reg[103][10] + loc_oh_reg[104][10] + loc_oh_reg[105][10] + loc_oh_reg[106][10] + loc_oh_reg[107][10] + loc_oh_reg[108][10] + loc_oh_reg[109][10] + loc_oh_reg[110][10] + loc_oh_reg[111][10] + loc_oh_reg[112][10] + loc_oh_reg[113][10] + loc_oh_reg[114][10] + loc_oh_reg[115][10] + loc_oh_reg[116][10] + loc_oh_reg[117][10] + loc_oh_reg[118][10] + loc_oh_reg[119][10] + loc_oh_reg[120][10] + loc_oh_reg[121][10] + loc_oh_reg[122][10] + loc_oh_reg[123][10] + loc_oh_reg[124][10] + loc_oh_reg[125][10] + loc_oh_reg[126][10] + loc_oh_reg[127][10];
    n_dsum_reg[84] = loc_oh_reg[128][10] + loc_oh_reg[129][10] + loc_oh_reg[130][10] + loc_oh_reg[131][10] + loc_oh_reg[132][10] + loc_oh_reg[133][10] + loc_oh_reg[134][10] + loc_oh_reg[135][10] + loc_oh_reg[136][10] + loc_oh_reg[137][10] + loc_oh_reg[138][10] + loc_oh_reg[139][10] + loc_oh_reg[140][10] + loc_oh_reg[141][10] + loc_oh_reg[142][10] + loc_oh_reg[143][10] + loc_oh_reg[144][10] + loc_oh_reg[145][10] + loc_oh_reg[146][10] + loc_oh_reg[147][10] + loc_oh_reg[148][10] + loc_oh_reg[149][10] + loc_oh_reg[150][10] + loc_oh_reg[151][10] + loc_oh_reg[152][10] + loc_oh_reg[153][10] + loc_oh_reg[154][10] + loc_oh_reg[155][10] + loc_oh_reg[156][10] + loc_oh_reg[157][10] + loc_oh_reg[158][10] + loc_oh_reg[159][10];
    n_dsum_reg[85] = loc_oh_reg[160][10] + loc_oh_reg[161][10] + loc_oh_reg[162][10] + loc_oh_reg[163][10] + loc_oh_reg[164][10] + loc_oh_reg[165][10] + loc_oh_reg[166][10] + loc_oh_reg[167][10] + loc_oh_reg[168][10] + loc_oh_reg[169][10] + loc_oh_reg[170][10] + loc_oh_reg[171][10] + loc_oh_reg[172][10] + loc_oh_reg[173][10] + loc_oh_reg[174][10] + loc_oh_reg[175][10] + loc_oh_reg[176][10] + loc_oh_reg[177][10] + loc_oh_reg[178][10] + loc_oh_reg[179][10] + loc_oh_reg[180][10] + loc_oh_reg[181][10] + loc_oh_reg[182][10] + loc_oh_reg[183][10] + loc_oh_reg[184][10] + loc_oh_reg[185][10] + loc_oh_reg[186][10] + loc_oh_reg[187][10] + loc_oh_reg[188][10] + loc_oh_reg[189][10] + loc_oh_reg[190][10] + loc_oh_reg[191][10];
    n_dsum_reg[86] = loc_oh_reg[192][10] + loc_oh_reg[193][10] + loc_oh_reg[194][10] + loc_oh_reg[195][10] + loc_oh_reg[196][10] + loc_oh_reg[197][10] + loc_oh_reg[198][10] + loc_oh_reg[199][10] + loc_oh_reg[200][10] + loc_oh_reg[201][10] + loc_oh_reg[202][10] + loc_oh_reg[203][10] + loc_oh_reg[204][10] + loc_oh_reg[205][10] + loc_oh_reg[206][10] + loc_oh_reg[207][10] + loc_oh_reg[208][10] + loc_oh_reg[209][10] + loc_oh_reg[210][10] + loc_oh_reg[211][10] + loc_oh_reg[212][10] + loc_oh_reg[213][10] + loc_oh_reg[214][10] + loc_oh_reg[215][10] + loc_oh_reg[216][10] + loc_oh_reg[217][10] + loc_oh_reg[218][10] + loc_oh_reg[219][10] + loc_oh_reg[220][10] + loc_oh_reg[221][10] + loc_oh_reg[222][10] + loc_oh_reg[223][10];
    n_dsum_reg[87] = loc_oh_reg[224][10] + loc_oh_reg[225][10] + loc_oh_reg[226][10] + loc_oh_reg[227][10] + loc_oh_reg[228][10] + loc_oh_reg[229][10] + loc_oh_reg[230][10] + loc_oh_reg[231][10] + loc_oh_reg[232][10] + loc_oh_reg[233][10] + loc_oh_reg[234][10] + loc_oh_reg[235][10] + loc_oh_reg[236][10] + loc_oh_reg[237][10] + loc_oh_reg[238][10] + loc_oh_reg[239][10] + loc_oh_reg[240][10] + loc_oh_reg[241][10] + loc_oh_reg[242][10] + loc_oh_reg[243][10] + loc_oh_reg[244][10] + loc_oh_reg[245][10] + loc_oh_reg[246][10] + loc_oh_reg[247][10] + loc_oh_reg[248][10] + loc_oh_reg[249][10] + loc_oh_reg[250][10] + loc_oh_reg[251][10] + loc_oh_reg[252][10] + loc_oh_reg[253][10] + loc_oh_reg[254][10] + loc_oh_reg[255][10];

    n_dsum_reg[88] = loc_oh_reg[0][11] + loc_oh_reg[1][11] + loc_oh_reg[2][11] + loc_oh_reg[3][11] + loc_oh_reg[4][11] + loc_oh_reg[5][11] + loc_oh_reg[6][11] + loc_oh_reg[7][11] + loc_oh_reg[8][11] + loc_oh_reg[9][11] + loc_oh_reg[10][11] + loc_oh_reg[11][11] + loc_oh_reg[12][11] + loc_oh_reg[13][11] + loc_oh_reg[14][11] + loc_oh_reg[15][11] + loc_oh_reg[16][11] + loc_oh_reg[17][11] + loc_oh_reg[18][11] + loc_oh_reg[19][11] + loc_oh_reg[20][11] + loc_oh_reg[21][11] + loc_oh_reg[22][11] + loc_oh_reg[23][11] + loc_oh_reg[24][11] + loc_oh_reg[25][11] + loc_oh_reg[26][11] + loc_oh_reg[27][11] + loc_oh_reg[28][11] + loc_oh_reg[29][11] + loc_oh_reg[30][11] + loc_oh_reg[31][11];
    n_dsum_reg[89] = loc_oh_reg[32][11] + loc_oh_reg[33][11] + loc_oh_reg[34][11] + loc_oh_reg[35][11] + loc_oh_reg[36][11] + loc_oh_reg[37][11] + loc_oh_reg[38][11] + loc_oh_reg[39][11] + loc_oh_reg[40][11] + loc_oh_reg[41][11] + loc_oh_reg[42][11] + loc_oh_reg[43][11] + loc_oh_reg[44][11] + loc_oh_reg[45][11] + loc_oh_reg[46][11] + loc_oh_reg[47][11] + loc_oh_reg[48][11] + loc_oh_reg[49][11] + loc_oh_reg[50][11] + loc_oh_reg[51][11] + loc_oh_reg[52][11] + loc_oh_reg[53][11] + loc_oh_reg[54][11] + loc_oh_reg[55][11] + loc_oh_reg[56][11] + loc_oh_reg[57][11] + loc_oh_reg[58][11] + loc_oh_reg[59][11] + loc_oh_reg[60][11] + loc_oh_reg[61][11] + loc_oh_reg[62][11] + loc_oh_reg[63][11];
    n_dsum_reg[90] = loc_oh_reg[64][11] + loc_oh_reg[65][11] + loc_oh_reg[66][11] + loc_oh_reg[67][11] + loc_oh_reg[68][11] + loc_oh_reg[69][11] + loc_oh_reg[70][11] + loc_oh_reg[71][11] + loc_oh_reg[72][11] + loc_oh_reg[73][11] + loc_oh_reg[74][11] + loc_oh_reg[75][11] + loc_oh_reg[76][11] + loc_oh_reg[77][11] + loc_oh_reg[78][11] + loc_oh_reg[79][11] + loc_oh_reg[80][11] + loc_oh_reg[81][11] + loc_oh_reg[82][11] + loc_oh_reg[83][11] + loc_oh_reg[84][11] + loc_oh_reg[85][11] + loc_oh_reg[86][11] + loc_oh_reg[87][11] + loc_oh_reg[88][11] + loc_oh_reg[89][11] + loc_oh_reg[90][11] + loc_oh_reg[91][11] + loc_oh_reg[92][11] + loc_oh_reg[93][11] + loc_oh_reg[94][11] + loc_oh_reg[95][11];
    n_dsum_reg[91] = loc_oh_reg[96][11] + loc_oh_reg[97][11] + loc_oh_reg[98][11] + loc_oh_reg[99][11] + loc_oh_reg[100][11] + loc_oh_reg[101][11] + loc_oh_reg[102][11] + loc_oh_reg[103][11] + loc_oh_reg[104][11] + loc_oh_reg[105][11] + loc_oh_reg[106][11] + loc_oh_reg[107][11] + loc_oh_reg[108][11] + loc_oh_reg[109][11] + loc_oh_reg[110][11] + loc_oh_reg[111][11] + loc_oh_reg[112][11] + loc_oh_reg[113][11] + loc_oh_reg[114][11] + loc_oh_reg[115][11] + loc_oh_reg[116][11] + loc_oh_reg[117][11] + loc_oh_reg[118][11] + loc_oh_reg[119][11] + loc_oh_reg[120][11] + loc_oh_reg[121][11] + loc_oh_reg[122][11] + loc_oh_reg[123][11] + loc_oh_reg[124][11] + loc_oh_reg[125][11] + loc_oh_reg[126][11] + loc_oh_reg[127][11];
    n_dsum_reg[92] = loc_oh_reg[128][11] + loc_oh_reg[129][11] + loc_oh_reg[130][11] + loc_oh_reg[131][11] + loc_oh_reg[132][11] + loc_oh_reg[133][11] + loc_oh_reg[134][11] + loc_oh_reg[135][11] + loc_oh_reg[136][11] + loc_oh_reg[137][11] + loc_oh_reg[138][11] + loc_oh_reg[139][11] + loc_oh_reg[140][11] + loc_oh_reg[141][11] + loc_oh_reg[142][11] + loc_oh_reg[143][11] + loc_oh_reg[144][11] + loc_oh_reg[145][11] + loc_oh_reg[146][11] + loc_oh_reg[147][11] + loc_oh_reg[148][11] + loc_oh_reg[149][11] + loc_oh_reg[150][11] + loc_oh_reg[151][11] + loc_oh_reg[152][11] + loc_oh_reg[153][11] + loc_oh_reg[154][11] + loc_oh_reg[155][11] + loc_oh_reg[156][11] + loc_oh_reg[157][11] + loc_oh_reg[158][11] + loc_oh_reg[159][11];
    n_dsum_reg[93] = loc_oh_reg[160][11] + loc_oh_reg[161][11] + loc_oh_reg[162][11] + loc_oh_reg[163][11] + loc_oh_reg[164][11] + loc_oh_reg[165][11] + loc_oh_reg[166][11] + loc_oh_reg[167][11] + loc_oh_reg[168][11] + loc_oh_reg[169][11] + loc_oh_reg[170][11] + loc_oh_reg[171][11] + loc_oh_reg[172][11] + loc_oh_reg[173][11] + loc_oh_reg[174][11] + loc_oh_reg[175][11] + loc_oh_reg[176][11] + loc_oh_reg[177][11] + loc_oh_reg[178][11] + loc_oh_reg[179][11] + loc_oh_reg[180][11] + loc_oh_reg[181][11] + loc_oh_reg[182][11] + loc_oh_reg[183][11] + loc_oh_reg[184][11] + loc_oh_reg[185][11] + loc_oh_reg[186][11] + loc_oh_reg[187][11] + loc_oh_reg[188][11] + loc_oh_reg[189][11] + loc_oh_reg[190][11] + loc_oh_reg[191][11];
    n_dsum_reg[94] = loc_oh_reg[192][11] + loc_oh_reg[193][11] + loc_oh_reg[194][11] + loc_oh_reg[195][11] + loc_oh_reg[196][11] + loc_oh_reg[197][11] + loc_oh_reg[198][11] + loc_oh_reg[199][11] + loc_oh_reg[200][11] + loc_oh_reg[201][11] + loc_oh_reg[202][11] + loc_oh_reg[203][11] + loc_oh_reg[204][11] + loc_oh_reg[205][11] + loc_oh_reg[206][11] + loc_oh_reg[207][11] + loc_oh_reg[208][11] + loc_oh_reg[209][11] + loc_oh_reg[210][11] + loc_oh_reg[211][11] + loc_oh_reg[212][11] + loc_oh_reg[213][11] + loc_oh_reg[214][11] + loc_oh_reg[215][11] + loc_oh_reg[216][11] + loc_oh_reg[217][11] + loc_oh_reg[218][11] + loc_oh_reg[219][11] + loc_oh_reg[220][11] + loc_oh_reg[221][11] + loc_oh_reg[222][11] + loc_oh_reg[223][11];
    n_dsum_reg[95] = loc_oh_reg[224][11] + loc_oh_reg[225][11] + loc_oh_reg[226][11] + loc_oh_reg[227][11] + loc_oh_reg[228][11] + loc_oh_reg[229][11] + loc_oh_reg[230][11] + loc_oh_reg[231][11] + loc_oh_reg[232][11] + loc_oh_reg[233][11] + loc_oh_reg[234][11] + loc_oh_reg[235][11] + loc_oh_reg[236][11] + loc_oh_reg[237][11] + loc_oh_reg[238][11] + loc_oh_reg[239][11] + loc_oh_reg[240][11] + loc_oh_reg[241][11] + loc_oh_reg[242][11] + loc_oh_reg[243][11] + loc_oh_reg[244][11] + loc_oh_reg[245][11] + loc_oh_reg[246][11] + loc_oh_reg[247][11] + loc_oh_reg[248][11] + loc_oh_reg[249][11] + loc_oh_reg[250][11] + loc_oh_reg[251][11] + loc_oh_reg[252][11] + loc_oh_reg[253][11] + loc_oh_reg[254][11] + loc_oh_reg[255][11];

    n_dsum_reg[96] = loc_oh_reg[0][12] + loc_oh_reg[1][12] + loc_oh_reg[2][12] + loc_oh_reg[3][12] + loc_oh_reg[4][12] + loc_oh_reg[5][12] + loc_oh_reg[6][12] + loc_oh_reg[7][12] + loc_oh_reg[8][12] + loc_oh_reg[9][12] + loc_oh_reg[10][12] + loc_oh_reg[11][12] + loc_oh_reg[12][12] + loc_oh_reg[13][12] + loc_oh_reg[14][12] + loc_oh_reg[15][12] + loc_oh_reg[16][12] + loc_oh_reg[17][12] + loc_oh_reg[18][12] + loc_oh_reg[19][12] + loc_oh_reg[20][12] + loc_oh_reg[21][12] + loc_oh_reg[22][12] + loc_oh_reg[23][12] + loc_oh_reg[24][12] + loc_oh_reg[25][12] + loc_oh_reg[26][12] + loc_oh_reg[27][12] + loc_oh_reg[28][12] + loc_oh_reg[29][12] + loc_oh_reg[30][12] + loc_oh_reg[31][12];
    n_dsum_reg[97] = loc_oh_reg[32][12] + loc_oh_reg[33][12] + loc_oh_reg[34][12] + loc_oh_reg[35][12] + loc_oh_reg[36][12] + loc_oh_reg[37][12] + loc_oh_reg[38][12] + loc_oh_reg[39][12] + loc_oh_reg[40][12] + loc_oh_reg[41][12] + loc_oh_reg[42][12] + loc_oh_reg[43][12] + loc_oh_reg[44][12] + loc_oh_reg[45][12] + loc_oh_reg[46][12] + loc_oh_reg[47][12] + loc_oh_reg[48][12] + loc_oh_reg[49][12] + loc_oh_reg[50][12] + loc_oh_reg[51][12] + loc_oh_reg[52][12] + loc_oh_reg[53][12] + loc_oh_reg[54][12] + loc_oh_reg[55][12] + loc_oh_reg[56][12] + loc_oh_reg[57][12] + loc_oh_reg[58][12] + loc_oh_reg[59][12] + loc_oh_reg[60][12] + loc_oh_reg[61][12] + loc_oh_reg[62][12] + loc_oh_reg[63][12];
    n_dsum_reg[98] = loc_oh_reg[64][12] + loc_oh_reg[65][12] + loc_oh_reg[66][12] + loc_oh_reg[67][12] + loc_oh_reg[68][12] + loc_oh_reg[69][12] + loc_oh_reg[70][12] + loc_oh_reg[71][12] + loc_oh_reg[72][12] + loc_oh_reg[73][12] + loc_oh_reg[74][12] + loc_oh_reg[75][12] + loc_oh_reg[76][12] + loc_oh_reg[77][12] + loc_oh_reg[78][12] + loc_oh_reg[79][12] + loc_oh_reg[80][12] + loc_oh_reg[81][12] + loc_oh_reg[82][12] + loc_oh_reg[83][12] + loc_oh_reg[84][12] + loc_oh_reg[85][12] + loc_oh_reg[86][12] + loc_oh_reg[87][12] + loc_oh_reg[88][12] + loc_oh_reg[89][12] + loc_oh_reg[90][12] + loc_oh_reg[91][12] + loc_oh_reg[92][12] + loc_oh_reg[93][12] + loc_oh_reg[94][12] + loc_oh_reg[95][12];
    n_dsum_reg[99] = loc_oh_reg[96][12] + loc_oh_reg[97][12] + loc_oh_reg[98][12] + loc_oh_reg[99][12] + loc_oh_reg[100][12] + loc_oh_reg[101][12] + loc_oh_reg[102][12] + loc_oh_reg[103][12] + loc_oh_reg[104][12] + loc_oh_reg[105][12] + loc_oh_reg[106][12] + loc_oh_reg[107][12] + loc_oh_reg[108][12] + loc_oh_reg[109][12] + loc_oh_reg[110][12] + loc_oh_reg[111][12] + loc_oh_reg[112][12] + loc_oh_reg[113][12] + loc_oh_reg[114][12] + loc_oh_reg[115][12] + loc_oh_reg[116][12] + loc_oh_reg[117][12] + loc_oh_reg[118][12] + loc_oh_reg[119][12] + loc_oh_reg[120][12] + loc_oh_reg[121][12] + loc_oh_reg[122][12] + loc_oh_reg[123][12] + loc_oh_reg[124][12] + loc_oh_reg[125][12] + loc_oh_reg[126][12] + loc_oh_reg[127][12];
    n_dsum_reg[100] = loc_oh_reg[128][12] + loc_oh_reg[129][12] + loc_oh_reg[130][12] + loc_oh_reg[131][12] + loc_oh_reg[132][12] + loc_oh_reg[133][12] + loc_oh_reg[134][12] + loc_oh_reg[135][12] + loc_oh_reg[136][12] + loc_oh_reg[137][12] + loc_oh_reg[138][12] + loc_oh_reg[139][12] + loc_oh_reg[140][12] + loc_oh_reg[141][12] + loc_oh_reg[142][12] + loc_oh_reg[143][12] + loc_oh_reg[144][12] + loc_oh_reg[145][12] + loc_oh_reg[146][12] + loc_oh_reg[147][12] + loc_oh_reg[148][12] + loc_oh_reg[149][12] + loc_oh_reg[150][12] + loc_oh_reg[151][12] + loc_oh_reg[152][12] + loc_oh_reg[153][12] + loc_oh_reg[154][12] + loc_oh_reg[155][12] + loc_oh_reg[156][12] + loc_oh_reg[157][12] + loc_oh_reg[158][12] + loc_oh_reg[159][12];
    n_dsum_reg[101] = loc_oh_reg[160][12] + loc_oh_reg[161][12] + loc_oh_reg[162][12] + loc_oh_reg[163][12] + loc_oh_reg[164][12] + loc_oh_reg[165][12] + loc_oh_reg[166][12] + loc_oh_reg[167][12] + loc_oh_reg[168][12] + loc_oh_reg[169][12] + loc_oh_reg[170][12] + loc_oh_reg[171][12] + loc_oh_reg[172][12] + loc_oh_reg[173][12] + loc_oh_reg[174][12] + loc_oh_reg[175][12] + loc_oh_reg[176][12] + loc_oh_reg[177][12] + loc_oh_reg[178][12] + loc_oh_reg[179][12] + loc_oh_reg[180][12] + loc_oh_reg[181][12] + loc_oh_reg[182][12] + loc_oh_reg[183][12] + loc_oh_reg[184][12] + loc_oh_reg[185][12] + loc_oh_reg[186][12] + loc_oh_reg[187][12] + loc_oh_reg[188][12] + loc_oh_reg[189][12] + loc_oh_reg[190][12] + loc_oh_reg[191][12];
    n_dsum_reg[102] = loc_oh_reg[192][12] + loc_oh_reg[193][12] + loc_oh_reg[194][12] + loc_oh_reg[195][12] + loc_oh_reg[196][12] + loc_oh_reg[197][12] + loc_oh_reg[198][12] + loc_oh_reg[199][12] + loc_oh_reg[200][12] + loc_oh_reg[201][12] + loc_oh_reg[202][12] + loc_oh_reg[203][12] + loc_oh_reg[204][12] + loc_oh_reg[205][12] + loc_oh_reg[206][12] + loc_oh_reg[207][12] + loc_oh_reg[208][12] + loc_oh_reg[209][12] + loc_oh_reg[210][12] + loc_oh_reg[211][12] + loc_oh_reg[212][12] + loc_oh_reg[213][12] + loc_oh_reg[214][12] + loc_oh_reg[215][12] + loc_oh_reg[216][12] + loc_oh_reg[217][12] + loc_oh_reg[218][12] + loc_oh_reg[219][12] + loc_oh_reg[220][12] + loc_oh_reg[221][12] + loc_oh_reg[222][12] + loc_oh_reg[223][12];
    n_dsum_reg[103] = loc_oh_reg[224][12] + loc_oh_reg[225][12] + loc_oh_reg[226][12] + loc_oh_reg[227][12] + loc_oh_reg[228][12] + loc_oh_reg[229][12] + loc_oh_reg[230][12] + loc_oh_reg[231][12] + loc_oh_reg[232][12] + loc_oh_reg[233][12] + loc_oh_reg[234][12] + loc_oh_reg[235][12] + loc_oh_reg[236][12] + loc_oh_reg[237][12] + loc_oh_reg[238][12] + loc_oh_reg[239][12] + loc_oh_reg[240][12] + loc_oh_reg[241][12] + loc_oh_reg[242][12] + loc_oh_reg[243][12] + loc_oh_reg[244][12] + loc_oh_reg[245][12] + loc_oh_reg[246][12] + loc_oh_reg[247][12] + loc_oh_reg[248][12] + loc_oh_reg[249][12] + loc_oh_reg[250][12] + loc_oh_reg[251][12] + loc_oh_reg[252][12] + loc_oh_reg[253][12] + loc_oh_reg[254][12] + loc_oh_reg[255][12];

    n_dsum_reg[104] = loc_oh_reg[0][13] + loc_oh_reg[1][13] + loc_oh_reg[2][13] + loc_oh_reg[3][13] + loc_oh_reg[4][13] + loc_oh_reg[5][13] + loc_oh_reg[6][13] + loc_oh_reg[7][13] + loc_oh_reg[8][13] + loc_oh_reg[9][13] + loc_oh_reg[10][13] + loc_oh_reg[11][13] + loc_oh_reg[12][13] + loc_oh_reg[13][13] + loc_oh_reg[14][13] + loc_oh_reg[15][13] + loc_oh_reg[16][13] + loc_oh_reg[17][13] + loc_oh_reg[18][13] + loc_oh_reg[19][13] + loc_oh_reg[20][13] + loc_oh_reg[21][13] + loc_oh_reg[22][13] + loc_oh_reg[23][13] + loc_oh_reg[24][13] + loc_oh_reg[25][13] + loc_oh_reg[26][13] + loc_oh_reg[27][13] + loc_oh_reg[28][13] + loc_oh_reg[29][13] + loc_oh_reg[30][13] + loc_oh_reg[31][13];
    n_dsum_reg[105] = loc_oh_reg[32][13] + loc_oh_reg[33][13] + loc_oh_reg[34][13] + loc_oh_reg[35][13] + loc_oh_reg[36][13] + loc_oh_reg[37][13] + loc_oh_reg[38][13] + loc_oh_reg[39][13] + loc_oh_reg[40][13] + loc_oh_reg[41][13] + loc_oh_reg[42][13] + loc_oh_reg[43][13] + loc_oh_reg[44][13] + loc_oh_reg[45][13] + loc_oh_reg[46][13] + loc_oh_reg[47][13] + loc_oh_reg[48][13] + loc_oh_reg[49][13] + loc_oh_reg[50][13] + loc_oh_reg[51][13] + loc_oh_reg[52][13] + loc_oh_reg[53][13] + loc_oh_reg[54][13] + loc_oh_reg[55][13] + loc_oh_reg[56][13] + loc_oh_reg[57][13] + loc_oh_reg[58][13] + loc_oh_reg[59][13] + loc_oh_reg[60][13] + loc_oh_reg[61][13] + loc_oh_reg[62][13] + loc_oh_reg[63][13];
    n_dsum_reg[106] = loc_oh_reg[64][13] + loc_oh_reg[65][13] + loc_oh_reg[66][13] + loc_oh_reg[67][13] + loc_oh_reg[68][13] + loc_oh_reg[69][13] + loc_oh_reg[70][13] + loc_oh_reg[71][13] + loc_oh_reg[72][13] + loc_oh_reg[73][13] + loc_oh_reg[74][13] + loc_oh_reg[75][13] + loc_oh_reg[76][13] + loc_oh_reg[77][13] + loc_oh_reg[78][13] + loc_oh_reg[79][13] + loc_oh_reg[80][13] + loc_oh_reg[81][13] + loc_oh_reg[82][13] + loc_oh_reg[83][13] + loc_oh_reg[84][13] + loc_oh_reg[85][13] + loc_oh_reg[86][13] + loc_oh_reg[87][13] + loc_oh_reg[88][13] + loc_oh_reg[89][13] + loc_oh_reg[90][13] + loc_oh_reg[91][13] + loc_oh_reg[92][13] + loc_oh_reg[93][13] + loc_oh_reg[94][13] + loc_oh_reg[95][13];
    n_dsum_reg[107] = loc_oh_reg[96][13] + loc_oh_reg[97][13] + loc_oh_reg[98][13] + loc_oh_reg[99][13] + loc_oh_reg[100][13] + loc_oh_reg[101][13] + loc_oh_reg[102][13] + loc_oh_reg[103][13] + loc_oh_reg[104][13] + loc_oh_reg[105][13] + loc_oh_reg[106][13] + loc_oh_reg[107][13] + loc_oh_reg[108][13] + loc_oh_reg[109][13] + loc_oh_reg[110][13] + loc_oh_reg[111][13] + loc_oh_reg[112][13] + loc_oh_reg[113][13] + loc_oh_reg[114][13] + loc_oh_reg[115][13] + loc_oh_reg[116][13] + loc_oh_reg[117][13] + loc_oh_reg[118][13] + loc_oh_reg[119][13] + loc_oh_reg[120][13] + loc_oh_reg[121][13] + loc_oh_reg[122][13] + loc_oh_reg[123][13] + loc_oh_reg[124][13] + loc_oh_reg[125][13] + loc_oh_reg[126][13] + loc_oh_reg[127][13];
    n_dsum_reg[108] = loc_oh_reg[128][13] + loc_oh_reg[129][13] + loc_oh_reg[130][13] + loc_oh_reg[131][13] + loc_oh_reg[132][13] + loc_oh_reg[133][13] + loc_oh_reg[134][13] + loc_oh_reg[135][13] + loc_oh_reg[136][13] + loc_oh_reg[137][13] + loc_oh_reg[138][13] + loc_oh_reg[139][13] + loc_oh_reg[140][13] + loc_oh_reg[141][13] + loc_oh_reg[142][13] + loc_oh_reg[143][13] + loc_oh_reg[144][13] + loc_oh_reg[145][13] + loc_oh_reg[146][13] + loc_oh_reg[147][13] + loc_oh_reg[148][13] + loc_oh_reg[149][13] + loc_oh_reg[150][13] + loc_oh_reg[151][13] + loc_oh_reg[152][13] + loc_oh_reg[153][13] + loc_oh_reg[154][13] + loc_oh_reg[155][13] + loc_oh_reg[156][13] + loc_oh_reg[157][13] + loc_oh_reg[158][13] + loc_oh_reg[159][13];
    n_dsum_reg[109] = loc_oh_reg[160][13] + loc_oh_reg[161][13] + loc_oh_reg[162][13] + loc_oh_reg[163][13] + loc_oh_reg[164][13] + loc_oh_reg[165][13] + loc_oh_reg[166][13] + loc_oh_reg[167][13] + loc_oh_reg[168][13] + loc_oh_reg[169][13] + loc_oh_reg[170][13] + loc_oh_reg[171][13] + loc_oh_reg[172][13] + loc_oh_reg[173][13] + loc_oh_reg[174][13] + loc_oh_reg[175][13] + loc_oh_reg[176][13] + loc_oh_reg[177][13] + loc_oh_reg[178][13] + loc_oh_reg[179][13] + loc_oh_reg[180][13] + loc_oh_reg[181][13] + loc_oh_reg[182][13] + loc_oh_reg[183][13] + loc_oh_reg[184][13] + loc_oh_reg[185][13] + loc_oh_reg[186][13] + loc_oh_reg[187][13] + loc_oh_reg[188][13] + loc_oh_reg[189][13] + loc_oh_reg[190][13] + loc_oh_reg[191][13];
    n_dsum_reg[110] = loc_oh_reg[192][13] + loc_oh_reg[193][13] + loc_oh_reg[194][13] + loc_oh_reg[195][13] + loc_oh_reg[196][13] + loc_oh_reg[197][13] + loc_oh_reg[198][13] + loc_oh_reg[199][13] + loc_oh_reg[200][13] + loc_oh_reg[201][13] + loc_oh_reg[202][13] + loc_oh_reg[203][13] + loc_oh_reg[204][13] + loc_oh_reg[205][13] + loc_oh_reg[206][13] + loc_oh_reg[207][13] + loc_oh_reg[208][13] + loc_oh_reg[209][13] + loc_oh_reg[210][13] + loc_oh_reg[211][13] + loc_oh_reg[212][13] + loc_oh_reg[213][13] + loc_oh_reg[214][13] + loc_oh_reg[215][13] + loc_oh_reg[216][13] + loc_oh_reg[217][13] + loc_oh_reg[218][13] + loc_oh_reg[219][13] + loc_oh_reg[220][13] + loc_oh_reg[221][13] + loc_oh_reg[222][13] + loc_oh_reg[223][13];
    n_dsum_reg[111] = loc_oh_reg[224][13] + loc_oh_reg[225][13] + loc_oh_reg[226][13] + loc_oh_reg[227][13] + loc_oh_reg[228][13] + loc_oh_reg[229][13] + loc_oh_reg[230][13] + loc_oh_reg[231][13] + loc_oh_reg[232][13] + loc_oh_reg[233][13] + loc_oh_reg[234][13] + loc_oh_reg[235][13] + loc_oh_reg[236][13] + loc_oh_reg[237][13] + loc_oh_reg[238][13] + loc_oh_reg[239][13] + loc_oh_reg[240][13] + loc_oh_reg[241][13] + loc_oh_reg[242][13] + loc_oh_reg[243][13] + loc_oh_reg[244][13] + loc_oh_reg[245][13] + loc_oh_reg[246][13] + loc_oh_reg[247][13] + loc_oh_reg[248][13] + loc_oh_reg[249][13] + loc_oh_reg[250][13] + loc_oh_reg[251][13] + loc_oh_reg[252][13] + loc_oh_reg[253][13] + loc_oh_reg[254][13] + loc_oh_reg[255][13];

    n_dsum_reg[112] = loc_oh_reg[0][14] + loc_oh_reg[1][14] + loc_oh_reg[2][14] + loc_oh_reg[3][14] + loc_oh_reg[4][14] + loc_oh_reg[5][14] + loc_oh_reg[6][14] + loc_oh_reg[7][14] + loc_oh_reg[8][14] + loc_oh_reg[9][14] + loc_oh_reg[10][14] + loc_oh_reg[11][14] + loc_oh_reg[12][14] + loc_oh_reg[13][14] + loc_oh_reg[14][14] + loc_oh_reg[15][14] + loc_oh_reg[16][14] + loc_oh_reg[17][14] + loc_oh_reg[18][14] + loc_oh_reg[19][14] + loc_oh_reg[20][14] + loc_oh_reg[21][14] + loc_oh_reg[22][14] + loc_oh_reg[23][14] + loc_oh_reg[24][14] + loc_oh_reg[25][14] + loc_oh_reg[26][14] + loc_oh_reg[27][14] + loc_oh_reg[28][14] + loc_oh_reg[29][14] + loc_oh_reg[30][14] + loc_oh_reg[31][14];
    n_dsum_reg[113] = loc_oh_reg[32][14] + loc_oh_reg[33][14] + loc_oh_reg[34][14] + loc_oh_reg[35][14] + loc_oh_reg[36][14] + loc_oh_reg[37][14] + loc_oh_reg[38][14] + loc_oh_reg[39][14] + loc_oh_reg[40][14] + loc_oh_reg[41][14] + loc_oh_reg[42][14] + loc_oh_reg[43][14] + loc_oh_reg[44][14] + loc_oh_reg[45][14] + loc_oh_reg[46][14] + loc_oh_reg[47][14] + loc_oh_reg[48][14] + loc_oh_reg[49][14] + loc_oh_reg[50][14] + loc_oh_reg[51][14] + loc_oh_reg[52][14] + loc_oh_reg[53][14] + loc_oh_reg[54][14] + loc_oh_reg[55][14] + loc_oh_reg[56][14] + loc_oh_reg[57][14] + loc_oh_reg[58][14] + loc_oh_reg[59][14] + loc_oh_reg[60][14] + loc_oh_reg[61][14] + loc_oh_reg[62][14] + loc_oh_reg[63][14];
    n_dsum_reg[114] = loc_oh_reg[64][14] + loc_oh_reg[65][14] + loc_oh_reg[66][14] + loc_oh_reg[67][14] + loc_oh_reg[68][14] + loc_oh_reg[69][14] + loc_oh_reg[70][14] + loc_oh_reg[71][14] + loc_oh_reg[72][14] + loc_oh_reg[73][14] + loc_oh_reg[74][14] + loc_oh_reg[75][14] + loc_oh_reg[76][14] + loc_oh_reg[77][14] + loc_oh_reg[78][14] + loc_oh_reg[79][14] + loc_oh_reg[80][14] + loc_oh_reg[81][14] + loc_oh_reg[82][14] + loc_oh_reg[83][14] + loc_oh_reg[84][14] + loc_oh_reg[85][14] + loc_oh_reg[86][14] + loc_oh_reg[87][14] + loc_oh_reg[88][14] + loc_oh_reg[89][14] + loc_oh_reg[90][14] + loc_oh_reg[91][14] + loc_oh_reg[92][14] + loc_oh_reg[93][14] + loc_oh_reg[94][14] + loc_oh_reg[95][14];
    n_dsum_reg[115] = loc_oh_reg[96][14] + loc_oh_reg[97][14] + loc_oh_reg[98][14] + loc_oh_reg[99][14] + loc_oh_reg[100][14] + loc_oh_reg[101][14] + loc_oh_reg[102][14] + loc_oh_reg[103][14] + loc_oh_reg[104][14] + loc_oh_reg[105][14] + loc_oh_reg[106][14] + loc_oh_reg[107][14] + loc_oh_reg[108][14] + loc_oh_reg[109][14] + loc_oh_reg[110][14] + loc_oh_reg[111][14] + loc_oh_reg[112][14] + loc_oh_reg[113][14] + loc_oh_reg[114][14] + loc_oh_reg[115][14] + loc_oh_reg[116][14] + loc_oh_reg[117][14] + loc_oh_reg[118][14] + loc_oh_reg[119][14] + loc_oh_reg[120][14] + loc_oh_reg[121][14] + loc_oh_reg[122][14] + loc_oh_reg[123][14] + loc_oh_reg[124][14] + loc_oh_reg[125][14] + loc_oh_reg[126][14] + loc_oh_reg[127][14];
    n_dsum_reg[116] = loc_oh_reg[128][14] + loc_oh_reg[129][14] + loc_oh_reg[130][14] + loc_oh_reg[131][14] + loc_oh_reg[132][14] + loc_oh_reg[133][14] + loc_oh_reg[134][14] + loc_oh_reg[135][14] + loc_oh_reg[136][14] + loc_oh_reg[137][14] + loc_oh_reg[138][14] + loc_oh_reg[139][14] + loc_oh_reg[140][14] + loc_oh_reg[141][14] + loc_oh_reg[142][14] + loc_oh_reg[143][14] + loc_oh_reg[144][14] + loc_oh_reg[145][14] + loc_oh_reg[146][14] + loc_oh_reg[147][14] + loc_oh_reg[148][14] + loc_oh_reg[149][14] + loc_oh_reg[150][14] + loc_oh_reg[151][14] + loc_oh_reg[152][14] + loc_oh_reg[153][14] + loc_oh_reg[154][14] + loc_oh_reg[155][14] + loc_oh_reg[156][14] + loc_oh_reg[157][14] + loc_oh_reg[158][14] + loc_oh_reg[159][14];
    n_dsum_reg[117] = loc_oh_reg[160][14] + loc_oh_reg[161][14] + loc_oh_reg[162][14] + loc_oh_reg[163][14] + loc_oh_reg[164][14] + loc_oh_reg[165][14] + loc_oh_reg[166][14] + loc_oh_reg[167][14] + loc_oh_reg[168][14] + loc_oh_reg[169][14] + loc_oh_reg[170][14] + loc_oh_reg[171][14] + loc_oh_reg[172][14] + loc_oh_reg[173][14] + loc_oh_reg[174][14] + loc_oh_reg[175][14] + loc_oh_reg[176][14] + loc_oh_reg[177][14] + loc_oh_reg[178][14] + loc_oh_reg[179][14] + loc_oh_reg[180][14] + loc_oh_reg[181][14] + loc_oh_reg[182][14] + loc_oh_reg[183][14] + loc_oh_reg[184][14] + loc_oh_reg[185][14] + loc_oh_reg[186][14] + loc_oh_reg[187][14] + loc_oh_reg[188][14] + loc_oh_reg[189][14] + loc_oh_reg[190][14] + loc_oh_reg[191][14];
    n_dsum_reg[118] = loc_oh_reg[192][14] + loc_oh_reg[193][14] + loc_oh_reg[194][14] + loc_oh_reg[195][14] + loc_oh_reg[196][14] + loc_oh_reg[197][14] + loc_oh_reg[198][14] + loc_oh_reg[199][14] + loc_oh_reg[200][14] + loc_oh_reg[201][14] + loc_oh_reg[202][14] + loc_oh_reg[203][14] + loc_oh_reg[204][14] + loc_oh_reg[205][14] + loc_oh_reg[206][14] + loc_oh_reg[207][14] + loc_oh_reg[208][14] + loc_oh_reg[209][14] + loc_oh_reg[210][14] + loc_oh_reg[211][14] + loc_oh_reg[212][14] + loc_oh_reg[213][14] + loc_oh_reg[214][14] + loc_oh_reg[215][14] + loc_oh_reg[216][14] + loc_oh_reg[217][14] + loc_oh_reg[218][14] + loc_oh_reg[219][14] + loc_oh_reg[220][14] + loc_oh_reg[221][14] + loc_oh_reg[222][14] + loc_oh_reg[223][14];
    n_dsum_reg[119] = loc_oh_reg[224][14] + loc_oh_reg[225][14] + loc_oh_reg[226][14] + loc_oh_reg[227][14] + loc_oh_reg[228][14] + loc_oh_reg[229][14] + loc_oh_reg[230][14] + loc_oh_reg[231][14] + loc_oh_reg[232][14] + loc_oh_reg[233][14] + loc_oh_reg[234][14] + loc_oh_reg[235][14] + loc_oh_reg[236][14] + loc_oh_reg[237][14] + loc_oh_reg[238][14] + loc_oh_reg[239][14] + loc_oh_reg[240][14] + loc_oh_reg[241][14] + loc_oh_reg[242][14] + loc_oh_reg[243][14] + loc_oh_reg[244][14] + loc_oh_reg[245][14] + loc_oh_reg[246][14] + loc_oh_reg[247][14] + loc_oh_reg[248][14] + loc_oh_reg[249][14] + loc_oh_reg[250][14] + loc_oh_reg[251][14] + loc_oh_reg[252][14] + loc_oh_reg[253][14] + loc_oh_reg[254][14] + loc_oh_reg[255][14];

    n_dsum_reg[120] = loc_oh_reg[0][15] + loc_oh_reg[1][15] + loc_oh_reg[2][15] + loc_oh_reg[3][15] + loc_oh_reg[4][15] + loc_oh_reg[5][15] + loc_oh_reg[6][15] + loc_oh_reg[7][15] + loc_oh_reg[8][15] + loc_oh_reg[9][15] + loc_oh_reg[10][15] + loc_oh_reg[11][15] + loc_oh_reg[12][15] + loc_oh_reg[13][15] + loc_oh_reg[14][15] + loc_oh_reg[15][15] + loc_oh_reg[16][15] + loc_oh_reg[17][15] + loc_oh_reg[18][15] + loc_oh_reg[19][15] + loc_oh_reg[20][15] + loc_oh_reg[21][15] + loc_oh_reg[22][15] + loc_oh_reg[23][15] + loc_oh_reg[24][15] + loc_oh_reg[25][15] + loc_oh_reg[26][15] + loc_oh_reg[27][15] + loc_oh_reg[28][15] + loc_oh_reg[29][15] + loc_oh_reg[30][15] + loc_oh_reg[31][15];
    n_dsum_reg[121] = loc_oh_reg[32][15] + loc_oh_reg[33][15] + loc_oh_reg[34][15] + loc_oh_reg[35][15] + loc_oh_reg[36][15] + loc_oh_reg[37][15] + loc_oh_reg[38][15] + loc_oh_reg[39][15] + loc_oh_reg[40][15] + loc_oh_reg[41][15] + loc_oh_reg[42][15] + loc_oh_reg[43][15] + loc_oh_reg[44][15] + loc_oh_reg[45][15] + loc_oh_reg[46][15] + loc_oh_reg[47][15] + loc_oh_reg[48][15] + loc_oh_reg[49][15] + loc_oh_reg[50][15] + loc_oh_reg[51][15] + loc_oh_reg[52][15] + loc_oh_reg[53][15] + loc_oh_reg[54][15] + loc_oh_reg[55][15] + loc_oh_reg[56][15] + loc_oh_reg[57][15] + loc_oh_reg[58][15] + loc_oh_reg[59][15] + loc_oh_reg[60][15] + loc_oh_reg[61][15] + loc_oh_reg[62][15] + loc_oh_reg[63][15];
    n_dsum_reg[122] = loc_oh_reg[64][15] + loc_oh_reg[65][15] + loc_oh_reg[66][15] + loc_oh_reg[67][15] + loc_oh_reg[68][15] + loc_oh_reg[69][15] + loc_oh_reg[70][15] + loc_oh_reg[71][15] + loc_oh_reg[72][15] + loc_oh_reg[73][15] + loc_oh_reg[74][15] + loc_oh_reg[75][15] + loc_oh_reg[76][15] + loc_oh_reg[77][15] + loc_oh_reg[78][15] + loc_oh_reg[79][15] + loc_oh_reg[80][15] + loc_oh_reg[81][15] + loc_oh_reg[82][15] + loc_oh_reg[83][15] + loc_oh_reg[84][15] + loc_oh_reg[85][15] + loc_oh_reg[86][15] + loc_oh_reg[87][15] + loc_oh_reg[88][15] + loc_oh_reg[89][15] + loc_oh_reg[90][15] + loc_oh_reg[91][15] + loc_oh_reg[92][15] + loc_oh_reg[93][15] + loc_oh_reg[94][15] + loc_oh_reg[95][15];
    n_dsum_reg[123] = loc_oh_reg[96][15] + loc_oh_reg[97][15] + loc_oh_reg[98][15] + loc_oh_reg[99][15] + loc_oh_reg[100][15] + loc_oh_reg[101][15] + loc_oh_reg[102][15] + loc_oh_reg[103][15] + loc_oh_reg[104][15] + loc_oh_reg[105][15] + loc_oh_reg[106][15] + loc_oh_reg[107][15] + loc_oh_reg[108][15] + loc_oh_reg[109][15] + loc_oh_reg[110][15] + loc_oh_reg[111][15] + loc_oh_reg[112][15] + loc_oh_reg[113][15] + loc_oh_reg[114][15] + loc_oh_reg[115][15] + loc_oh_reg[116][15] + loc_oh_reg[117][15] + loc_oh_reg[118][15] + loc_oh_reg[119][15] + loc_oh_reg[120][15] + loc_oh_reg[121][15] + loc_oh_reg[122][15] + loc_oh_reg[123][15] + loc_oh_reg[124][15] + loc_oh_reg[125][15] + loc_oh_reg[126][15] + loc_oh_reg[127][15];
    n_dsum_reg[124] = loc_oh_reg[128][15] + loc_oh_reg[129][15] + loc_oh_reg[130][15] + loc_oh_reg[131][15] + loc_oh_reg[132][15] + loc_oh_reg[133][15] + loc_oh_reg[134][15] + loc_oh_reg[135][15] + loc_oh_reg[136][15] + loc_oh_reg[137][15] + loc_oh_reg[138][15] + loc_oh_reg[139][15] + loc_oh_reg[140][15] + loc_oh_reg[141][15] + loc_oh_reg[142][15] + loc_oh_reg[143][15] + loc_oh_reg[144][15] + loc_oh_reg[145][15] + loc_oh_reg[146][15] + loc_oh_reg[147][15] + loc_oh_reg[148][15] + loc_oh_reg[149][15] + loc_oh_reg[150][15] + loc_oh_reg[151][15] + loc_oh_reg[152][15] + loc_oh_reg[153][15] + loc_oh_reg[154][15] + loc_oh_reg[155][15] + loc_oh_reg[156][15] + loc_oh_reg[157][15] + loc_oh_reg[158][15] + loc_oh_reg[159][15];
    n_dsum_reg[125] = loc_oh_reg[160][15] + loc_oh_reg[161][15] + loc_oh_reg[162][15] + loc_oh_reg[163][15] + loc_oh_reg[164][15] + loc_oh_reg[165][15] + loc_oh_reg[166][15] + loc_oh_reg[167][15] + loc_oh_reg[168][15] + loc_oh_reg[169][15] + loc_oh_reg[170][15] + loc_oh_reg[171][15] + loc_oh_reg[172][15] + loc_oh_reg[173][15] + loc_oh_reg[174][15] + loc_oh_reg[175][15] + loc_oh_reg[176][15] + loc_oh_reg[177][15] + loc_oh_reg[178][15] + loc_oh_reg[179][15] + loc_oh_reg[180][15] + loc_oh_reg[181][15] + loc_oh_reg[182][15] + loc_oh_reg[183][15] + loc_oh_reg[184][15] + loc_oh_reg[185][15] + loc_oh_reg[186][15] + loc_oh_reg[187][15] + loc_oh_reg[188][15] + loc_oh_reg[189][15] + loc_oh_reg[190][15] + loc_oh_reg[191][15];
    n_dsum_reg[126] = loc_oh_reg[192][15] + loc_oh_reg[193][15] + loc_oh_reg[194][15] + loc_oh_reg[195][15] + loc_oh_reg[196][15] + loc_oh_reg[197][15] + loc_oh_reg[198][15] + loc_oh_reg[199][15] + loc_oh_reg[200][15] + loc_oh_reg[201][15] + loc_oh_reg[202][15] + loc_oh_reg[203][15] + loc_oh_reg[204][15] + loc_oh_reg[205][15] + loc_oh_reg[206][15] + loc_oh_reg[207][15] + loc_oh_reg[208][15] + loc_oh_reg[209][15] + loc_oh_reg[210][15] + loc_oh_reg[211][15] + loc_oh_reg[212][15] + loc_oh_reg[213][15] + loc_oh_reg[214][15] + loc_oh_reg[215][15] + loc_oh_reg[216][15] + loc_oh_reg[217][15] + loc_oh_reg[218][15] + loc_oh_reg[219][15] + loc_oh_reg[220][15] + loc_oh_reg[221][15] + loc_oh_reg[222][15] + loc_oh_reg[223][15];
    n_dsum_reg[127] = loc_oh_reg[224][15] + loc_oh_reg[225][15] + loc_oh_reg[226][15] + loc_oh_reg[227][15] + loc_oh_reg[228][15] + loc_oh_reg[229][15] + loc_oh_reg[230][15] + loc_oh_reg[231][15] + loc_oh_reg[232][15] + loc_oh_reg[233][15] + loc_oh_reg[234][15] + loc_oh_reg[235][15] + loc_oh_reg[236][15] + loc_oh_reg[237][15] + loc_oh_reg[238][15] + loc_oh_reg[239][15] + loc_oh_reg[240][15] + loc_oh_reg[241][15] + loc_oh_reg[242][15] + loc_oh_reg[243][15] + loc_oh_reg[244][15] + loc_oh_reg[245][15] + loc_oh_reg[246][15] + loc_oh_reg[247][15] + loc_oh_reg[248][15] + loc_oh_reg[249][15] + loc_oh_reg[250][15] + loc_oh_reg[251][15] + loc_oh_reg[252][15] + loc_oh_reg[253][15] + loc_oh_reg[254][15] + loc_oh_reg[255][15];
end

// COMB3: get part_reg
always@* begin
    if(part_en) begin
        n_part_reg[0] = dsum_reg[0] + dsum_reg[1] + dsum_reg[2] + dsum_reg[3] + dsum_reg[4] + dsum_reg[5] + dsum_reg[6] + dsum_reg[7];
        n_part_reg[1] = dsum_reg[8] + dsum_reg[9] + dsum_reg[10] + dsum_reg[11] + dsum_reg[12] + dsum_reg[13] + dsum_reg[14] + dsum_reg[15];
        n_part_reg[2] = dsum_reg[16] + dsum_reg[17] + dsum_reg[18] + dsum_reg[19] + dsum_reg[20] + dsum_reg[21] + dsum_reg[22] + dsum_reg[23];
        n_part_reg[3] = dsum_reg[24] + dsum_reg[25] + dsum_reg[26] + dsum_reg[27] + dsum_reg[28] + dsum_reg[29] + dsum_reg[30] + dsum_reg[31];
        n_part_reg[4] = dsum_reg[32] + dsum_reg[33] + dsum_reg[34] + dsum_reg[35] + dsum_reg[36] + dsum_reg[37] + dsum_reg[38] + dsum_reg[39];
        n_part_reg[5] = dsum_reg[40] + dsum_reg[41] + dsum_reg[42] + dsum_reg[43] + dsum_reg[44] + dsum_reg[45] + dsum_reg[46] + dsum_reg[47];
        n_part_reg[6] = dsum_reg[48] + dsum_reg[49] + dsum_reg[50] + dsum_reg[51] + dsum_reg[52] + dsum_reg[53] + dsum_reg[54] + dsum_reg[55];
        n_part_reg[7] = dsum_reg[56] + dsum_reg[57] + dsum_reg[58] + dsum_reg[59] + dsum_reg[60] + dsum_reg[61] + dsum_reg[62] + dsum_reg[63];
        n_part_reg[8] = dsum_reg[64] + dsum_reg[65] + dsum_reg[66] + dsum_reg[67] + dsum_reg[68] + dsum_reg[69] + dsum_reg[70] + dsum_reg[71];
        n_part_reg[9] = dsum_reg[72] + dsum_reg[73] + dsum_reg[74] + dsum_reg[75] + dsum_reg[76] + dsum_reg[77] + dsum_reg[78] + dsum_reg[79];
        n_part_reg[10] = dsum_reg[80] + dsum_reg[81] + dsum_reg[82] + dsum_reg[83] + dsum_reg[84] + dsum_reg[85] + dsum_reg[86] + dsum_reg[87];
        n_part_reg[11] = dsum_reg[88] + dsum_reg[89] + dsum_reg[90] + dsum_reg[91] + dsum_reg[92] + dsum_reg[93] + dsum_reg[94] + dsum_reg[95];
        n_part_reg[12] = dsum_reg[96] + dsum_reg[97] + dsum_reg[98] + dsum_reg[99] + dsum_reg[100] + dsum_reg[101] + dsum_reg[102] + dsum_reg[103];
        n_part_reg[13] = dsum_reg[104] + dsum_reg[105] + dsum_reg[106] + dsum_reg[107] + dsum_reg[108] + dsum_reg[109] + dsum_reg[110] + dsum_reg[111];
        n_part_reg[14] = dsum_reg[112] + dsum_reg[113] + dsum_reg[114] + dsum_reg[115] + dsum_reg[116] + dsum_reg[117] + dsum_reg[118] + dsum_reg[119];
        n_part_reg[15] = dsum_reg[120] + dsum_reg[121] + dsum_reg[122] + dsum_reg[123] + dsum_reg[124] + dsum_reg[125] + dsum_reg[126] + dsum_reg[127];
    end else begin
        n_part_reg[0] = part_reg[0] + dsum_reg[0] + dsum_reg[1] + dsum_reg[2] + dsum_reg[3] + dsum_reg[4] + dsum_reg[5] + dsum_reg[6] + dsum_reg[7];
        n_part_reg[1] = part_reg[1] + dsum_reg[8] + dsum_reg[9] + dsum_reg[10] + dsum_reg[11] + dsum_reg[12] + dsum_reg[13] + dsum_reg[14] + dsum_reg[15];
        n_part_reg[2] = part_reg[2] + dsum_reg[16] + dsum_reg[17] + dsum_reg[18] + dsum_reg[19] + dsum_reg[20] + dsum_reg[21] + dsum_reg[22] + dsum_reg[23];
        n_part_reg[3] = part_reg[3] + dsum_reg[24] + dsum_reg[25] + dsum_reg[26] + dsum_reg[27] + dsum_reg[28] + dsum_reg[29] + dsum_reg[30] + dsum_reg[31];
        n_part_reg[4] = part_reg[4] + dsum_reg[32] + dsum_reg[33] + dsum_reg[34] + dsum_reg[35] + dsum_reg[36] + dsum_reg[37] + dsum_reg[38] + dsum_reg[39];
        n_part_reg[5] = part_reg[5] + dsum_reg[40] + dsum_reg[41] + dsum_reg[42] + dsum_reg[43] + dsum_reg[44] + dsum_reg[45] + dsum_reg[46] + dsum_reg[47];
        n_part_reg[6] = part_reg[6] + dsum_reg[48] + dsum_reg[49] + dsum_reg[50] + dsum_reg[51] + dsum_reg[52] + dsum_reg[53] + dsum_reg[54] + dsum_reg[55];
        n_part_reg[7] = part_reg[7] + dsum_reg[56] + dsum_reg[57] + dsum_reg[58] + dsum_reg[59] + dsum_reg[60] + dsum_reg[61] + dsum_reg[62] + dsum_reg[63];
        n_part_reg[8] = part_reg[8] + dsum_reg[64] + dsum_reg[65] + dsum_reg[66] + dsum_reg[67] + dsum_reg[68] + dsum_reg[69] + dsum_reg[70] + dsum_reg[71];
        n_part_reg[9] = part_reg[9] + dsum_reg[72] + dsum_reg[73] + dsum_reg[74] + dsum_reg[75] + dsum_reg[76] + dsum_reg[77] + dsum_reg[78] + dsum_reg[79];
        n_part_reg[10] = part_reg[10] + dsum_reg[80] + dsum_reg[81] + dsum_reg[82] + dsum_reg[83] + dsum_reg[84] + dsum_reg[85] + dsum_reg[86] + dsum_reg[87];
        n_part_reg[11] = part_reg[11] + dsum_reg[88] + dsum_reg[89] + dsum_reg[90] + dsum_reg[91] + dsum_reg[92] + dsum_reg[93] + dsum_reg[94] + dsum_reg[95];
        n_part_reg[12] = part_reg[12] + dsum_reg[96] + dsum_reg[97] + dsum_reg[98] + dsum_reg[99] + dsum_reg[100] + dsum_reg[101] + dsum_reg[102] + dsum_reg[103];
        n_part_reg[13] = part_reg[13] + dsum_reg[104] + dsum_reg[105] + dsum_reg[106] + dsum_reg[107] + dsum_reg[108] + dsum_reg[109] + dsum_reg[110] + dsum_reg[111];
        n_part_reg[14] = part_reg[14] + dsum_reg[112] + dsum_reg[113] + dsum_reg[114] + dsum_reg[115] + dsum_reg[116] + dsum_reg[117] + dsum_reg[118] + dsum_reg[119];
        n_part_reg[15] = part_reg[15] + dsum_reg[120] + dsum_reg[121] + dsum_reg[122] + dsum_reg[123] + dsum_reg[124] + dsum_reg[125] + dsum_reg[126] + dsum_reg[127];
    end
end

// COMB4: comparator so as to get next
always@* begin
    // for work 0
    res0_comp[0] = (part_reg[1] >= part_reg[0]) ? {part_reg[1], 4'd1} : {part_reg[0], 4'd0};
    res0_comp[1] = (part_reg[2] >= part_reg[3]) ? {part_reg[2], 4'd2} : {part_reg[3], 4'd3};
    res0_comp[2] = (part_reg[4] >= part_reg[5]) ? {part_reg[4], 4'd4} : {part_reg[5], 4'd5};
    res0_comp[3] = (part_reg[6] >= part_reg[7]) ? {part_reg[6], 4'd6} : {part_reg[7], 4'd7};
    res0_comp[4] = (part_reg[8] >= part_reg[9]) ? {part_reg[8], 4'd8} : {part_reg[9], 4'd9};
    res0_comp[5] = (part_reg[10] >= part_reg[11]) ? {part_reg[10], 4'd10} : {part_reg[11], 4'd11};
    res0_comp[6] = (part_reg[12] >= part_reg[13]) ? {part_reg[12], 4'd12} : {part_reg[13], 4'd13};
    res0_comp[7] = (part_reg[14] >= part_reg[15]) ? {part_reg[14], 4'd14} : {part_reg[15], 4'd15};

    res1_comp[0] = (res0_comp[0][11:4] >= res0_comp[1][11:4]) ? res0_comp[0] : res0_comp[1];
    res1_comp[1] = (res0_comp[2][11:4] >= res0_comp[3][11:4]) ? res0_comp[2] : res0_comp[3];
    res1_comp[2] = (res0_comp[4][11:4] >= res0_comp[5][11:4]) ? res0_comp[4] : res0_comp[5];
    res1_comp[3] = (res0_comp[6][11:4] >= res0_comp[7][11:4]) ? res0_comp[6] : res0_comp[7];

    res2_comp[0] = (res1_comp[0][11:4] >= res1_comp[1][11:4]) ? res1_comp[0] : res1_comp[1];
    res2_comp[1] = (res1_comp[2][11:4] >= res1_comp[3][11:4]) ? res1_comp[2] : res1_comp[3];

    res3_comp = (res2_comp[0][11:4] >= res2_comp[1][11:4]) ? res2_comp[0] : res2_comp[1];
end

always@* begin
	case(batch_num_reg[3:0])
		4'd1: n_next_wdata = {60'd0, res4_comp};
		4'd2: n_next_wdata = {56'd0, res4_comp, 4'd0};
		4'd3: n_next_wdata = {52'd0, res4_comp, 8'd0};
		4'd4: n_next_wdata = {48'd0, res4_comp, 12'd0};
		4'd5: n_next_wdata = {44'd0, res4_comp, 16'd0};
		4'd6: n_next_wdata = {40'd0, res4_comp, 20'd0};
		4'd7: n_next_wdata = {36'd0, res4_comp, 24'd0};
		4'd8: n_next_wdata = {32'd0, res4_comp, 28'd0};
		4'd9: n_next_wdata = {28'd0, res4_comp, 32'd0};
		4'd10: n_next_wdata = {24'd0, res4_comp, 36'd0};
		4'd11: n_next_wdata = {20'd0, res4_comp, 40'd0};
		4'd12: n_next_wdata = {16'd0, res4_comp, 44'd0};
		4'd13: n_next_wdata = {12'd0, res4_comp, 48'd0};
		4'd14: n_next_wdata = {8'd0, res4_comp, 52'd0};
		4'd15: n_next_wdata = {4'd0, res4_comp, 56'd0};
		4'd0: n_next_wdata = {res4_comp, 60'd0};
		default: n_next_wdata = 64'd0;
	endcase
end

always@* begin
	if(part_en) begin
		case(batch_num_reg[3:0])
			4'd1: n_next_bytemask = 16'b1111_1111_1111_1110;
			4'd2: n_next_bytemask = 16'b1111_1111_1111_1101;
			4'd3: n_next_bytemask = 16'b1111_1111_1111_1011;
			4'd4: n_next_bytemask = 16'b1111_1111_1111_0111;
			4'd5: n_next_bytemask = 16'b1111_1111_1110_1111;
			4'd6: n_next_bytemask = 16'b1111_1111_1101_1111;
			4'd7: n_next_bytemask = 16'b1111_1111_1011_1111;
			4'd8: n_next_bytemask = 16'b1111_1111_0111_1111;
			4'd9: n_next_bytemask = 16'b1111_1110_1111_1111;
			4'd10: n_next_bytemask = 16'b1111_1101_1111_1111;
			4'd11: n_next_bytemask = 16'b1111_1011_1111_1111;
			4'd12: n_next_bytemask = 16'b1111_0111_1111_1111;
			4'd13: n_next_bytemask = 16'b1110_1111_1111_1111;
			4'd14: n_next_bytemask = 16'b1101_1111_1111_1111;
			4'd15: n_next_bytemask = 16'b1011_1111_1111_1111;
			4'd0: n_next_bytemask = 16'b0111_1111_1111_1111;
			default: n_next_bytemask = 16'b1111_1111_1111_1111;
		endcase
			n_next_waddr = (batch_num_reg - 1) / 16;
	end else begin
		n_next_bytemask = 16'b1111_1111_1111_1111;
		n_next_waddr = next_waddr;
	end
end

// COMB5 proposal_cnt
always@* begin
	if(part_en) begin
		for(i = 0; i < 16; i = i + 1) begin
			if(res4_comp == i) begin
				n_proposal_cnt[i] = proposal_cnt[i] + 1;
			end else begin
				n_proposal_cnt[i] = proposal_cnt[i];
			end
		end
	end else begin
		for(i = 0; i < 16; i = i + 1) begin
			n_proposal_cnt[i] = proposal_cnt[i];
		end
	end
end

always@* begin
	case(batch_num_reg[3:0])
		4'd1: n_pro_wdata = {120'd0, proposal_cnt[res4_comp]};
		4'd2: n_pro_wdata = {112'd0, proposal_cnt[res4_comp], 8'd0};
		4'd3: n_pro_wdata = {104'd0, proposal_cnt[res4_comp], 16'd0};
		4'd4: n_pro_wdata = {96'd0, proposal_cnt[res4_comp], 24'd0};
		4'd5: n_pro_wdata = {88'd0, proposal_cnt[res4_comp], 32'd0};
		4'd6: n_pro_wdata = {80'd0, proposal_cnt[res4_comp], 40'd0};
		4'd7: n_pro_wdata = {72'd0, proposal_cnt[res4_comp], 48'd0};
		4'd8: n_pro_wdata = {64'd0, proposal_cnt[res4_comp], 56'd0};
		4'd9: n_pro_wdata = {56'd0, proposal_cnt[res4_comp], 64'd0};
		4'd10: n_pro_wdata = {48'd0, proposal_cnt[res4_comp], 72'd0};
		4'd11: n_pro_wdata = {40'd0, proposal_cnt[res4_comp], 80'd0};
		4'd12: n_pro_wdata = {32'd0, proposal_cnt[res4_comp], 88'd0};
		4'd13: n_pro_wdata = {24'd0, proposal_cnt[res4_comp], 96'd0};
		4'd14: n_pro_wdata = {16'd0, proposal_cnt[res4_comp], 104'd0};
		4'd15: n_pro_wdata = {8'd0, proposal_cnt[res4_comp], 112'd0};
		4'd0: n_pro_wdata = {proposal_cnt[res4_comp], 120'd0};
		default: n_pro_wdata = 128'd0;
	endcase
end

always@* begin
	if(part_en) begin
		case(batch_num_reg[3:0])
			4'd1: n_pro_bytemask = 16'b1111_1111_1111_1110;
			4'd2: n_pro_bytemask = 16'b1111_1111_1111_1101;
			4'd3: n_pro_bytemask = 16'b1111_1111_1111_1011;
			4'd4: n_pro_bytemask = 16'b1111_1111_1111_0111;
			4'd5: n_pro_bytemask = 16'b1111_1111_1110_1111;
			4'd6: n_pro_bytemask = 16'b1111_1111_1101_1111;
			4'd7: n_pro_bytemask = 16'b1111_1111_1011_1111;
			4'd8: n_pro_bytemask = 16'b1111_1111_0111_1111;
			4'd9: n_pro_bytemask = 16'b1111_1110_1111_1111;
			4'd10: n_pro_bytemask = 16'b1111_1101_1111_1111;
			4'd11: n_pro_bytemask = 16'b1111_1011_1111_1111;
			4'd12: n_pro_bytemask = 16'b1111_0111_1111_1111;
			4'd13: n_pro_bytemask = 16'b1110_1111_1111_1111;
			4'd14: n_pro_bytemask = 16'b1101_1111_1111_1111;
			4'd15: n_pro_bytemask = 16'b1011_1111_1111_1111;
			4'd0: n_pro_bytemask = 16'b0111_1111_1111_1111;
			default: n_pro_bytemask = 16'b1111_1111_1111_1111;
		endcase
			n_pro_waddr = (batch_num_reg - 1) / 16;
	end else begin
		n_pro_bytemask = 16'b1111_1111_1111_1111;
		n_pro_waddr = pro_waddr;
	end
end

always@* begin
	if(part_en) n_wen = 1;
	else n_wen = 0;
end

// TEST_CYCLE 2.0 -> slack -0.56
// TEST_CYCLE 2.5 -> slack -0.0225
// TEST_CYCLE 2.6 -> slack -0.1021
// TEST_CYCLE 3.0 -> slack 0

endmodule